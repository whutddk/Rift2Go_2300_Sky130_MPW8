magic
tech sky130A
magscale 1 2
timestamp 1671597917
<< obsli1 >>
rect 1104 2159 356408 428145
<< obsm1 >>
rect 566 2128 357498 428324
<< metal2 >>
rect 6458 429996 6514 430796
rect 16302 429996 16358 430796
rect 26146 429996 26202 430796
rect 35990 429996 36046 430796
rect 45834 429996 45890 430796
rect 55678 429996 55734 430796
rect 65522 429996 65578 430796
rect 75366 429996 75422 430796
rect 85210 429996 85266 430796
rect 95054 429996 95110 430796
rect 104898 429996 104954 430796
rect 114742 429996 114798 430796
rect 124586 429996 124642 430796
rect 134430 429996 134486 430796
rect 144274 429996 144330 430796
rect 154118 429996 154174 430796
rect 163962 429996 164018 430796
rect 173806 429996 173862 430796
rect 183650 429996 183706 430796
rect 193494 429996 193550 430796
rect 203338 429996 203394 430796
rect 213182 429996 213238 430796
rect 223026 429996 223082 430796
rect 232870 429996 232926 430796
rect 242714 429996 242770 430796
rect 252558 429996 252614 430796
rect 262402 429996 262458 430796
rect 272246 429996 272302 430796
rect 282090 429996 282146 430796
rect 291934 429996 291990 430796
rect 301778 429996 301834 430796
rect 311622 429996 311678 430796
rect 321466 429996 321522 430796
rect 331310 429996 331366 430796
rect 341154 429996 341210 430796
rect 350998 429996 351054 430796
rect 19982 0 20038 800
rect 20626 0 20682 800
rect 21270 0 21326 800
rect 21914 0 21970 800
rect 22558 0 22614 800
rect 23202 0 23258 800
rect 23846 0 23902 800
rect 24490 0 24546 800
rect 25134 0 25190 800
rect 25778 0 25834 800
rect 26422 0 26478 800
rect 27066 0 27122 800
rect 27710 0 27766 800
rect 28354 0 28410 800
rect 28998 0 29054 800
rect 29642 0 29698 800
rect 30286 0 30342 800
rect 30930 0 30986 800
rect 31574 0 31630 800
rect 32218 0 32274 800
rect 32862 0 32918 800
rect 33506 0 33562 800
rect 34150 0 34206 800
rect 34794 0 34850 800
rect 35438 0 35494 800
rect 36082 0 36138 800
rect 36726 0 36782 800
rect 37370 0 37426 800
rect 38014 0 38070 800
rect 38658 0 38714 800
rect 39302 0 39358 800
rect 39946 0 40002 800
rect 40590 0 40646 800
rect 41234 0 41290 800
rect 41878 0 41934 800
rect 42522 0 42578 800
rect 43166 0 43222 800
rect 43810 0 43866 800
rect 44454 0 44510 800
rect 45098 0 45154 800
rect 45742 0 45798 800
rect 46386 0 46442 800
rect 47030 0 47086 800
rect 47674 0 47730 800
rect 48318 0 48374 800
rect 48962 0 49018 800
rect 49606 0 49662 800
rect 50250 0 50306 800
rect 50894 0 50950 800
rect 51538 0 51594 800
rect 52182 0 52238 800
rect 52826 0 52882 800
rect 53470 0 53526 800
rect 54114 0 54170 800
rect 54758 0 54814 800
rect 55402 0 55458 800
rect 56046 0 56102 800
rect 56690 0 56746 800
rect 57334 0 57390 800
rect 57978 0 58034 800
rect 58622 0 58678 800
rect 59266 0 59322 800
rect 59910 0 59966 800
rect 60554 0 60610 800
rect 61198 0 61254 800
rect 61842 0 61898 800
rect 62486 0 62542 800
rect 63130 0 63186 800
rect 63774 0 63830 800
rect 64418 0 64474 800
rect 65062 0 65118 800
rect 65706 0 65762 800
rect 66350 0 66406 800
rect 66994 0 67050 800
rect 67638 0 67694 800
rect 68282 0 68338 800
rect 68926 0 68982 800
rect 69570 0 69626 800
rect 70214 0 70270 800
rect 70858 0 70914 800
rect 71502 0 71558 800
rect 72146 0 72202 800
rect 72790 0 72846 800
rect 73434 0 73490 800
rect 74078 0 74134 800
rect 74722 0 74778 800
rect 75366 0 75422 800
rect 76010 0 76066 800
rect 76654 0 76710 800
rect 77298 0 77354 800
rect 77942 0 77998 800
rect 78586 0 78642 800
rect 79230 0 79286 800
rect 79874 0 79930 800
rect 80518 0 80574 800
rect 81162 0 81218 800
rect 81806 0 81862 800
rect 82450 0 82506 800
rect 83094 0 83150 800
rect 83738 0 83794 800
rect 84382 0 84438 800
rect 85026 0 85082 800
rect 85670 0 85726 800
rect 86314 0 86370 800
rect 86958 0 87014 800
rect 87602 0 87658 800
rect 88246 0 88302 800
rect 88890 0 88946 800
rect 89534 0 89590 800
rect 90178 0 90234 800
rect 90822 0 90878 800
rect 91466 0 91522 800
rect 92110 0 92166 800
rect 92754 0 92810 800
rect 93398 0 93454 800
rect 94042 0 94098 800
rect 94686 0 94742 800
rect 95330 0 95386 800
rect 95974 0 96030 800
rect 96618 0 96674 800
rect 97262 0 97318 800
rect 97906 0 97962 800
rect 98550 0 98606 800
rect 99194 0 99250 800
rect 99838 0 99894 800
rect 100482 0 100538 800
rect 101126 0 101182 800
rect 101770 0 101826 800
rect 102414 0 102470 800
rect 103058 0 103114 800
rect 103702 0 103758 800
rect 104346 0 104402 800
rect 104990 0 105046 800
rect 105634 0 105690 800
rect 106278 0 106334 800
rect 106922 0 106978 800
rect 107566 0 107622 800
rect 108210 0 108266 800
rect 108854 0 108910 800
rect 109498 0 109554 800
rect 110142 0 110198 800
rect 110786 0 110842 800
rect 111430 0 111486 800
rect 112074 0 112130 800
rect 112718 0 112774 800
rect 113362 0 113418 800
rect 114006 0 114062 800
rect 114650 0 114706 800
rect 115294 0 115350 800
rect 115938 0 115994 800
rect 116582 0 116638 800
rect 117226 0 117282 800
rect 117870 0 117926 800
rect 118514 0 118570 800
rect 119158 0 119214 800
rect 119802 0 119858 800
rect 120446 0 120502 800
rect 121090 0 121146 800
rect 121734 0 121790 800
rect 122378 0 122434 800
rect 123022 0 123078 800
rect 123666 0 123722 800
rect 124310 0 124366 800
rect 124954 0 125010 800
rect 125598 0 125654 800
rect 126242 0 126298 800
rect 126886 0 126942 800
rect 127530 0 127586 800
rect 128174 0 128230 800
rect 128818 0 128874 800
rect 129462 0 129518 800
rect 130106 0 130162 800
rect 130750 0 130806 800
rect 131394 0 131450 800
rect 132038 0 132094 800
rect 132682 0 132738 800
rect 133326 0 133382 800
rect 133970 0 134026 800
rect 134614 0 134670 800
rect 135258 0 135314 800
rect 135902 0 135958 800
rect 136546 0 136602 800
rect 137190 0 137246 800
rect 137834 0 137890 800
rect 138478 0 138534 800
rect 139122 0 139178 800
rect 139766 0 139822 800
rect 140410 0 140466 800
rect 141054 0 141110 800
rect 141698 0 141754 800
rect 142342 0 142398 800
rect 142986 0 143042 800
rect 143630 0 143686 800
rect 144274 0 144330 800
rect 144918 0 144974 800
rect 145562 0 145618 800
rect 146206 0 146262 800
rect 146850 0 146906 800
rect 147494 0 147550 800
rect 148138 0 148194 800
rect 148782 0 148838 800
rect 149426 0 149482 800
rect 150070 0 150126 800
rect 150714 0 150770 800
rect 151358 0 151414 800
rect 152002 0 152058 800
rect 152646 0 152702 800
rect 153290 0 153346 800
rect 153934 0 153990 800
rect 154578 0 154634 800
rect 155222 0 155278 800
rect 155866 0 155922 800
rect 156510 0 156566 800
rect 157154 0 157210 800
rect 157798 0 157854 800
rect 158442 0 158498 800
rect 159086 0 159142 800
rect 159730 0 159786 800
rect 160374 0 160430 800
rect 161018 0 161074 800
rect 161662 0 161718 800
rect 162306 0 162362 800
rect 162950 0 163006 800
rect 163594 0 163650 800
rect 164238 0 164294 800
rect 164882 0 164938 800
rect 165526 0 165582 800
rect 166170 0 166226 800
rect 166814 0 166870 800
rect 167458 0 167514 800
rect 168102 0 168158 800
rect 168746 0 168802 800
rect 169390 0 169446 800
rect 170034 0 170090 800
rect 170678 0 170734 800
rect 171322 0 171378 800
rect 171966 0 172022 800
rect 172610 0 172666 800
rect 173254 0 173310 800
rect 173898 0 173954 800
rect 174542 0 174598 800
rect 175186 0 175242 800
rect 175830 0 175886 800
rect 176474 0 176530 800
rect 177118 0 177174 800
rect 177762 0 177818 800
rect 178406 0 178462 800
rect 179050 0 179106 800
rect 179694 0 179750 800
rect 180338 0 180394 800
rect 180982 0 181038 800
rect 181626 0 181682 800
rect 182270 0 182326 800
rect 182914 0 182970 800
rect 183558 0 183614 800
rect 184202 0 184258 800
rect 184846 0 184902 800
rect 185490 0 185546 800
rect 186134 0 186190 800
rect 186778 0 186834 800
rect 187422 0 187478 800
rect 188066 0 188122 800
rect 188710 0 188766 800
rect 189354 0 189410 800
rect 189998 0 190054 800
rect 190642 0 190698 800
rect 191286 0 191342 800
rect 191930 0 191986 800
rect 192574 0 192630 800
rect 193218 0 193274 800
rect 193862 0 193918 800
rect 194506 0 194562 800
rect 195150 0 195206 800
rect 195794 0 195850 800
rect 196438 0 196494 800
rect 197082 0 197138 800
rect 197726 0 197782 800
rect 198370 0 198426 800
rect 199014 0 199070 800
rect 199658 0 199714 800
rect 200302 0 200358 800
rect 200946 0 201002 800
rect 201590 0 201646 800
rect 202234 0 202290 800
rect 202878 0 202934 800
rect 203522 0 203578 800
rect 204166 0 204222 800
rect 204810 0 204866 800
rect 205454 0 205510 800
rect 206098 0 206154 800
rect 206742 0 206798 800
rect 207386 0 207442 800
rect 208030 0 208086 800
rect 208674 0 208730 800
rect 209318 0 209374 800
rect 209962 0 210018 800
rect 210606 0 210662 800
rect 211250 0 211306 800
rect 211894 0 211950 800
rect 212538 0 212594 800
rect 213182 0 213238 800
rect 213826 0 213882 800
rect 214470 0 214526 800
rect 215114 0 215170 800
rect 215758 0 215814 800
rect 216402 0 216458 800
rect 217046 0 217102 800
rect 217690 0 217746 800
rect 218334 0 218390 800
rect 218978 0 219034 800
rect 219622 0 219678 800
rect 220266 0 220322 800
rect 220910 0 220966 800
rect 221554 0 221610 800
rect 222198 0 222254 800
rect 222842 0 222898 800
rect 223486 0 223542 800
rect 224130 0 224186 800
rect 224774 0 224830 800
rect 225418 0 225474 800
rect 226062 0 226118 800
rect 226706 0 226762 800
rect 227350 0 227406 800
rect 227994 0 228050 800
rect 228638 0 228694 800
rect 229282 0 229338 800
rect 229926 0 229982 800
rect 230570 0 230626 800
rect 231214 0 231270 800
rect 231858 0 231914 800
rect 232502 0 232558 800
rect 233146 0 233202 800
rect 233790 0 233846 800
rect 234434 0 234490 800
rect 235078 0 235134 800
rect 235722 0 235778 800
rect 236366 0 236422 800
rect 237010 0 237066 800
rect 237654 0 237710 800
rect 238298 0 238354 800
rect 238942 0 238998 800
rect 239586 0 239642 800
rect 240230 0 240286 800
rect 240874 0 240930 800
rect 241518 0 241574 800
rect 242162 0 242218 800
rect 242806 0 242862 800
rect 243450 0 243506 800
rect 244094 0 244150 800
rect 244738 0 244794 800
rect 245382 0 245438 800
rect 246026 0 246082 800
rect 246670 0 246726 800
rect 247314 0 247370 800
rect 247958 0 248014 800
rect 248602 0 248658 800
rect 249246 0 249302 800
rect 249890 0 249946 800
rect 250534 0 250590 800
rect 251178 0 251234 800
rect 251822 0 251878 800
rect 252466 0 252522 800
rect 253110 0 253166 800
rect 253754 0 253810 800
rect 254398 0 254454 800
rect 255042 0 255098 800
rect 255686 0 255742 800
rect 256330 0 256386 800
rect 256974 0 257030 800
rect 257618 0 257674 800
rect 258262 0 258318 800
rect 258906 0 258962 800
rect 259550 0 259606 800
rect 260194 0 260250 800
rect 260838 0 260894 800
rect 261482 0 261538 800
rect 262126 0 262182 800
rect 262770 0 262826 800
rect 263414 0 263470 800
rect 264058 0 264114 800
rect 264702 0 264758 800
rect 265346 0 265402 800
rect 265990 0 266046 800
rect 266634 0 266690 800
rect 267278 0 267334 800
rect 267922 0 267978 800
rect 268566 0 268622 800
rect 269210 0 269266 800
rect 269854 0 269910 800
rect 270498 0 270554 800
rect 271142 0 271198 800
rect 271786 0 271842 800
rect 272430 0 272486 800
rect 273074 0 273130 800
rect 273718 0 273774 800
rect 274362 0 274418 800
rect 275006 0 275062 800
rect 275650 0 275706 800
rect 276294 0 276350 800
rect 276938 0 276994 800
rect 277582 0 277638 800
rect 278226 0 278282 800
rect 278870 0 278926 800
rect 279514 0 279570 800
rect 280158 0 280214 800
rect 280802 0 280858 800
rect 281446 0 281502 800
rect 282090 0 282146 800
rect 282734 0 282790 800
rect 283378 0 283434 800
rect 284022 0 284078 800
rect 284666 0 284722 800
rect 285310 0 285366 800
rect 285954 0 286010 800
rect 286598 0 286654 800
rect 287242 0 287298 800
rect 287886 0 287942 800
rect 288530 0 288586 800
rect 289174 0 289230 800
rect 289818 0 289874 800
rect 290462 0 290518 800
rect 291106 0 291162 800
rect 291750 0 291806 800
rect 292394 0 292450 800
rect 293038 0 293094 800
rect 293682 0 293738 800
rect 294326 0 294382 800
rect 294970 0 295026 800
rect 295614 0 295670 800
rect 296258 0 296314 800
rect 296902 0 296958 800
rect 297546 0 297602 800
rect 298190 0 298246 800
rect 298834 0 298890 800
rect 299478 0 299534 800
rect 300122 0 300178 800
rect 300766 0 300822 800
rect 301410 0 301466 800
rect 302054 0 302110 800
rect 302698 0 302754 800
rect 303342 0 303398 800
rect 303986 0 304042 800
rect 304630 0 304686 800
rect 305274 0 305330 800
rect 305918 0 305974 800
rect 306562 0 306618 800
rect 307206 0 307262 800
rect 307850 0 307906 800
rect 308494 0 308550 800
rect 309138 0 309194 800
rect 309782 0 309838 800
rect 310426 0 310482 800
rect 311070 0 311126 800
rect 311714 0 311770 800
rect 312358 0 312414 800
rect 313002 0 313058 800
rect 313646 0 313702 800
rect 314290 0 314346 800
rect 314934 0 314990 800
rect 315578 0 315634 800
rect 316222 0 316278 800
rect 316866 0 316922 800
rect 317510 0 317566 800
rect 318154 0 318210 800
rect 318798 0 318854 800
rect 319442 0 319498 800
rect 320086 0 320142 800
rect 320730 0 320786 800
rect 321374 0 321430 800
rect 322018 0 322074 800
rect 322662 0 322718 800
rect 323306 0 323362 800
rect 323950 0 324006 800
rect 324594 0 324650 800
rect 325238 0 325294 800
rect 325882 0 325938 800
rect 326526 0 326582 800
rect 327170 0 327226 800
rect 327814 0 327870 800
rect 328458 0 328514 800
rect 329102 0 329158 800
rect 329746 0 329802 800
rect 330390 0 330446 800
rect 331034 0 331090 800
rect 331678 0 331734 800
rect 332322 0 332378 800
rect 332966 0 333022 800
rect 333610 0 333666 800
rect 334254 0 334310 800
rect 334898 0 334954 800
rect 335542 0 335598 800
rect 336186 0 336242 800
rect 336830 0 336886 800
rect 337474 0 337530 800
<< obsm2 >>
rect 572 429940 6402 430114
rect 6570 429940 16246 430114
rect 16414 429940 26090 430114
rect 26258 429940 35934 430114
rect 36102 429940 45778 430114
rect 45946 429940 55622 430114
rect 55790 429940 65466 430114
rect 65634 429940 75310 430114
rect 75478 429940 85154 430114
rect 85322 429940 94998 430114
rect 95166 429940 104842 430114
rect 105010 429940 114686 430114
rect 114854 429940 124530 430114
rect 124698 429940 134374 430114
rect 134542 429940 144218 430114
rect 144386 429940 154062 430114
rect 154230 429940 163906 430114
rect 164074 429940 173750 430114
rect 173918 429940 183594 430114
rect 183762 429940 193438 430114
rect 193606 429940 203282 430114
rect 203450 429940 213126 430114
rect 213294 429940 222970 430114
rect 223138 429940 232814 430114
rect 232982 429940 242658 430114
rect 242826 429940 252502 430114
rect 252670 429940 262346 430114
rect 262514 429940 272190 430114
rect 272358 429940 282034 430114
rect 282202 429940 291878 430114
rect 292046 429940 301722 430114
rect 301890 429940 311566 430114
rect 311734 429940 321410 430114
rect 321578 429940 331254 430114
rect 331422 429940 341098 430114
rect 341266 429940 350942 430114
rect 351110 429940 357492 430114
rect 572 856 357492 429940
rect 572 800 19926 856
rect 20094 800 20570 856
rect 20738 800 21214 856
rect 21382 800 21858 856
rect 22026 800 22502 856
rect 22670 800 23146 856
rect 23314 800 23790 856
rect 23958 800 24434 856
rect 24602 800 25078 856
rect 25246 800 25722 856
rect 25890 800 26366 856
rect 26534 800 27010 856
rect 27178 800 27654 856
rect 27822 800 28298 856
rect 28466 800 28942 856
rect 29110 800 29586 856
rect 29754 800 30230 856
rect 30398 800 30874 856
rect 31042 800 31518 856
rect 31686 800 32162 856
rect 32330 800 32806 856
rect 32974 800 33450 856
rect 33618 800 34094 856
rect 34262 800 34738 856
rect 34906 800 35382 856
rect 35550 800 36026 856
rect 36194 800 36670 856
rect 36838 800 37314 856
rect 37482 800 37958 856
rect 38126 800 38602 856
rect 38770 800 39246 856
rect 39414 800 39890 856
rect 40058 800 40534 856
rect 40702 800 41178 856
rect 41346 800 41822 856
rect 41990 800 42466 856
rect 42634 800 43110 856
rect 43278 800 43754 856
rect 43922 800 44398 856
rect 44566 800 45042 856
rect 45210 800 45686 856
rect 45854 800 46330 856
rect 46498 800 46974 856
rect 47142 800 47618 856
rect 47786 800 48262 856
rect 48430 800 48906 856
rect 49074 800 49550 856
rect 49718 800 50194 856
rect 50362 800 50838 856
rect 51006 800 51482 856
rect 51650 800 52126 856
rect 52294 800 52770 856
rect 52938 800 53414 856
rect 53582 800 54058 856
rect 54226 800 54702 856
rect 54870 800 55346 856
rect 55514 800 55990 856
rect 56158 800 56634 856
rect 56802 800 57278 856
rect 57446 800 57922 856
rect 58090 800 58566 856
rect 58734 800 59210 856
rect 59378 800 59854 856
rect 60022 800 60498 856
rect 60666 800 61142 856
rect 61310 800 61786 856
rect 61954 800 62430 856
rect 62598 800 63074 856
rect 63242 800 63718 856
rect 63886 800 64362 856
rect 64530 800 65006 856
rect 65174 800 65650 856
rect 65818 800 66294 856
rect 66462 800 66938 856
rect 67106 800 67582 856
rect 67750 800 68226 856
rect 68394 800 68870 856
rect 69038 800 69514 856
rect 69682 800 70158 856
rect 70326 800 70802 856
rect 70970 800 71446 856
rect 71614 800 72090 856
rect 72258 800 72734 856
rect 72902 800 73378 856
rect 73546 800 74022 856
rect 74190 800 74666 856
rect 74834 800 75310 856
rect 75478 800 75954 856
rect 76122 800 76598 856
rect 76766 800 77242 856
rect 77410 800 77886 856
rect 78054 800 78530 856
rect 78698 800 79174 856
rect 79342 800 79818 856
rect 79986 800 80462 856
rect 80630 800 81106 856
rect 81274 800 81750 856
rect 81918 800 82394 856
rect 82562 800 83038 856
rect 83206 800 83682 856
rect 83850 800 84326 856
rect 84494 800 84970 856
rect 85138 800 85614 856
rect 85782 800 86258 856
rect 86426 800 86902 856
rect 87070 800 87546 856
rect 87714 800 88190 856
rect 88358 800 88834 856
rect 89002 800 89478 856
rect 89646 800 90122 856
rect 90290 800 90766 856
rect 90934 800 91410 856
rect 91578 800 92054 856
rect 92222 800 92698 856
rect 92866 800 93342 856
rect 93510 800 93986 856
rect 94154 800 94630 856
rect 94798 800 95274 856
rect 95442 800 95918 856
rect 96086 800 96562 856
rect 96730 800 97206 856
rect 97374 800 97850 856
rect 98018 800 98494 856
rect 98662 800 99138 856
rect 99306 800 99782 856
rect 99950 800 100426 856
rect 100594 800 101070 856
rect 101238 800 101714 856
rect 101882 800 102358 856
rect 102526 800 103002 856
rect 103170 800 103646 856
rect 103814 800 104290 856
rect 104458 800 104934 856
rect 105102 800 105578 856
rect 105746 800 106222 856
rect 106390 800 106866 856
rect 107034 800 107510 856
rect 107678 800 108154 856
rect 108322 800 108798 856
rect 108966 800 109442 856
rect 109610 800 110086 856
rect 110254 800 110730 856
rect 110898 800 111374 856
rect 111542 800 112018 856
rect 112186 800 112662 856
rect 112830 800 113306 856
rect 113474 800 113950 856
rect 114118 800 114594 856
rect 114762 800 115238 856
rect 115406 800 115882 856
rect 116050 800 116526 856
rect 116694 800 117170 856
rect 117338 800 117814 856
rect 117982 800 118458 856
rect 118626 800 119102 856
rect 119270 800 119746 856
rect 119914 800 120390 856
rect 120558 800 121034 856
rect 121202 800 121678 856
rect 121846 800 122322 856
rect 122490 800 122966 856
rect 123134 800 123610 856
rect 123778 800 124254 856
rect 124422 800 124898 856
rect 125066 800 125542 856
rect 125710 800 126186 856
rect 126354 800 126830 856
rect 126998 800 127474 856
rect 127642 800 128118 856
rect 128286 800 128762 856
rect 128930 800 129406 856
rect 129574 800 130050 856
rect 130218 800 130694 856
rect 130862 800 131338 856
rect 131506 800 131982 856
rect 132150 800 132626 856
rect 132794 800 133270 856
rect 133438 800 133914 856
rect 134082 800 134558 856
rect 134726 800 135202 856
rect 135370 800 135846 856
rect 136014 800 136490 856
rect 136658 800 137134 856
rect 137302 800 137778 856
rect 137946 800 138422 856
rect 138590 800 139066 856
rect 139234 800 139710 856
rect 139878 800 140354 856
rect 140522 800 140998 856
rect 141166 800 141642 856
rect 141810 800 142286 856
rect 142454 800 142930 856
rect 143098 800 143574 856
rect 143742 800 144218 856
rect 144386 800 144862 856
rect 145030 800 145506 856
rect 145674 800 146150 856
rect 146318 800 146794 856
rect 146962 800 147438 856
rect 147606 800 148082 856
rect 148250 800 148726 856
rect 148894 800 149370 856
rect 149538 800 150014 856
rect 150182 800 150658 856
rect 150826 800 151302 856
rect 151470 800 151946 856
rect 152114 800 152590 856
rect 152758 800 153234 856
rect 153402 800 153878 856
rect 154046 800 154522 856
rect 154690 800 155166 856
rect 155334 800 155810 856
rect 155978 800 156454 856
rect 156622 800 157098 856
rect 157266 800 157742 856
rect 157910 800 158386 856
rect 158554 800 159030 856
rect 159198 800 159674 856
rect 159842 800 160318 856
rect 160486 800 160962 856
rect 161130 800 161606 856
rect 161774 800 162250 856
rect 162418 800 162894 856
rect 163062 800 163538 856
rect 163706 800 164182 856
rect 164350 800 164826 856
rect 164994 800 165470 856
rect 165638 800 166114 856
rect 166282 800 166758 856
rect 166926 800 167402 856
rect 167570 800 168046 856
rect 168214 800 168690 856
rect 168858 800 169334 856
rect 169502 800 169978 856
rect 170146 800 170622 856
rect 170790 800 171266 856
rect 171434 800 171910 856
rect 172078 800 172554 856
rect 172722 800 173198 856
rect 173366 800 173842 856
rect 174010 800 174486 856
rect 174654 800 175130 856
rect 175298 800 175774 856
rect 175942 800 176418 856
rect 176586 800 177062 856
rect 177230 800 177706 856
rect 177874 800 178350 856
rect 178518 800 178994 856
rect 179162 800 179638 856
rect 179806 800 180282 856
rect 180450 800 180926 856
rect 181094 800 181570 856
rect 181738 800 182214 856
rect 182382 800 182858 856
rect 183026 800 183502 856
rect 183670 800 184146 856
rect 184314 800 184790 856
rect 184958 800 185434 856
rect 185602 800 186078 856
rect 186246 800 186722 856
rect 186890 800 187366 856
rect 187534 800 188010 856
rect 188178 800 188654 856
rect 188822 800 189298 856
rect 189466 800 189942 856
rect 190110 800 190586 856
rect 190754 800 191230 856
rect 191398 800 191874 856
rect 192042 800 192518 856
rect 192686 800 193162 856
rect 193330 800 193806 856
rect 193974 800 194450 856
rect 194618 800 195094 856
rect 195262 800 195738 856
rect 195906 800 196382 856
rect 196550 800 197026 856
rect 197194 800 197670 856
rect 197838 800 198314 856
rect 198482 800 198958 856
rect 199126 800 199602 856
rect 199770 800 200246 856
rect 200414 800 200890 856
rect 201058 800 201534 856
rect 201702 800 202178 856
rect 202346 800 202822 856
rect 202990 800 203466 856
rect 203634 800 204110 856
rect 204278 800 204754 856
rect 204922 800 205398 856
rect 205566 800 206042 856
rect 206210 800 206686 856
rect 206854 800 207330 856
rect 207498 800 207974 856
rect 208142 800 208618 856
rect 208786 800 209262 856
rect 209430 800 209906 856
rect 210074 800 210550 856
rect 210718 800 211194 856
rect 211362 800 211838 856
rect 212006 800 212482 856
rect 212650 800 213126 856
rect 213294 800 213770 856
rect 213938 800 214414 856
rect 214582 800 215058 856
rect 215226 800 215702 856
rect 215870 800 216346 856
rect 216514 800 216990 856
rect 217158 800 217634 856
rect 217802 800 218278 856
rect 218446 800 218922 856
rect 219090 800 219566 856
rect 219734 800 220210 856
rect 220378 800 220854 856
rect 221022 800 221498 856
rect 221666 800 222142 856
rect 222310 800 222786 856
rect 222954 800 223430 856
rect 223598 800 224074 856
rect 224242 800 224718 856
rect 224886 800 225362 856
rect 225530 800 226006 856
rect 226174 800 226650 856
rect 226818 800 227294 856
rect 227462 800 227938 856
rect 228106 800 228582 856
rect 228750 800 229226 856
rect 229394 800 229870 856
rect 230038 800 230514 856
rect 230682 800 231158 856
rect 231326 800 231802 856
rect 231970 800 232446 856
rect 232614 800 233090 856
rect 233258 800 233734 856
rect 233902 800 234378 856
rect 234546 800 235022 856
rect 235190 800 235666 856
rect 235834 800 236310 856
rect 236478 800 236954 856
rect 237122 800 237598 856
rect 237766 800 238242 856
rect 238410 800 238886 856
rect 239054 800 239530 856
rect 239698 800 240174 856
rect 240342 800 240818 856
rect 240986 800 241462 856
rect 241630 800 242106 856
rect 242274 800 242750 856
rect 242918 800 243394 856
rect 243562 800 244038 856
rect 244206 800 244682 856
rect 244850 800 245326 856
rect 245494 800 245970 856
rect 246138 800 246614 856
rect 246782 800 247258 856
rect 247426 800 247902 856
rect 248070 800 248546 856
rect 248714 800 249190 856
rect 249358 800 249834 856
rect 250002 800 250478 856
rect 250646 800 251122 856
rect 251290 800 251766 856
rect 251934 800 252410 856
rect 252578 800 253054 856
rect 253222 800 253698 856
rect 253866 800 254342 856
rect 254510 800 254986 856
rect 255154 800 255630 856
rect 255798 800 256274 856
rect 256442 800 256918 856
rect 257086 800 257562 856
rect 257730 800 258206 856
rect 258374 800 258850 856
rect 259018 800 259494 856
rect 259662 800 260138 856
rect 260306 800 260782 856
rect 260950 800 261426 856
rect 261594 800 262070 856
rect 262238 800 262714 856
rect 262882 800 263358 856
rect 263526 800 264002 856
rect 264170 800 264646 856
rect 264814 800 265290 856
rect 265458 800 265934 856
rect 266102 800 266578 856
rect 266746 800 267222 856
rect 267390 800 267866 856
rect 268034 800 268510 856
rect 268678 800 269154 856
rect 269322 800 269798 856
rect 269966 800 270442 856
rect 270610 800 271086 856
rect 271254 800 271730 856
rect 271898 800 272374 856
rect 272542 800 273018 856
rect 273186 800 273662 856
rect 273830 800 274306 856
rect 274474 800 274950 856
rect 275118 800 275594 856
rect 275762 800 276238 856
rect 276406 800 276882 856
rect 277050 800 277526 856
rect 277694 800 278170 856
rect 278338 800 278814 856
rect 278982 800 279458 856
rect 279626 800 280102 856
rect 280270 800 280746 856
rect 280914 800 281390 856
rect 281558 800 282034 856
rect 282202 800 282678 856
rect 282846 800 283322 856
rect 283490 800 283966 856
rect 284134 800 284610 856
rect 284778 800 285254 856
rect 285422 800 285898 856
rect 286066 800 286542 856
rect 286710 800 287186 856
rect 287354 800 287830 856
rect 287998 800 288474 856
rect 288642 800 289118 856
rect 289286 800 289762 856
rect 289930 800 290406 856
rect 290574 800 291050 856
rect 291218 800 291694 856
rect 291862 800 292338 856
rect 292506 800 292982 856
rect 293150 800 293626 856
rect 293794 800 294270 856
rect 294438 800 294914 856
rect 295082 800 295558 856
rect 295726 800 296202 856
rect 296370 800 296846 856
rect 297014 800 297490 856
rect 297658 800 298134 856
rect 298302 800 298778 856
rect 298946 800 299422 856
rect 299590 800 300066 856
rect 300234 800 300710 856
rect 300878 800 301354 856
rect 301522 800 301998 856
rect 302166 800 302642 856
rect 302810 800 303286 856
rect 303454 800 303930 856
rect 304098 800 304574 856
rect 304742 800 305218 856
rect 305386 800 305862 856
rect 306030 800 306506 856
rect 306674 800 307150 856
rect 307318 800 307794 856
rect 307962 800 308438 856
rect 308606 800 309082 856
rect 309250 800 309726 856
rect 309894 800 310370 856
rect 310538 800 311014 856
rect 311182 800 311658 856
rect 311826 800 312302 856
rect 312470 800 312946 856
rect 313114 800 313590 856
rect 313758 800 314234 856
rect 314402 800 314878 856
rect 315046 800 315522 856
rect 315690 800 316166 856
rect 316334 800 316810 856
rect 316978 800 317454 856
rect 317622 800 318098 856
rect 318266 800 318742 856
rect 318910 800 319386 856
rect 319554 800 320030 856
rect 320198 800 320674 856
rect 320842 800 321318 856
rect 321486 800 321962 856
rect 322130 800 322606 856
rect 322774 800 323250 856
rect 323418 800 323894 856
rect 324062 800 324538 856
rect 324706 800 325182 856
rect 325350 800 325826 856
rect 325994 800 326470 856
rect 326638 800 327114 856
rect 327282 800 327758 856
rect 327926 800 328402 856
rect 328570 800 329046 856
rect 329214 800 329690 856
rect 329858 800 330334 856
rect 330502 800 330978 856
rect 331146 800 331622 856
rect 331790 800 332266 856
rect 332434 800 332910 856
rect 333078 800 333554 856
rect 333722 800 334198 856
rect 334366 800 334842 856
rect 335010 800 335486 856
rect 335654 800 336130 856
rect 336298 800 336774 856
rect 336942 800 337418 856
rect 337586 800 357492 856
<< metal3 >>
rect 0 424328 800 424448
rect 356778 423920 357578 424040
rect 0 416440 800 416560
rect 356778 415896 357578 416016
rect 0 408552 800 408672
rect 356778 407872 357578 407992
rect 0 400664 800 400784
rect 356778 399848 357578 399968
rect 0 392776 800 392896
rect 356778 391824 357578 391944
rect 0 384888 800 385008
rect 356778 383800 357578 383920
rect 0 377000 800 377120
rect 356778 375776 357578 375896
rect 0 369112 800 369232
rect 356778 367752 357578 367872
rect 0 361224 800 361344
rect 356778 359728 357578 359848
rect 0 353336 800 353456
rect 356778 351704 357578 351824
rect 0 345448 800 345568
rect 356778 343680 357578 343800
rect 0 337560 800 337680
rect 356778 335656 357578 335776
rect 0 329672 800 329792
rect 356778 327632 357578 327752
rect 0 321784 800 321904
rect 356778 319608 357578 319728
rect 0 313896 800 314016
rect 356778 311584 357578 311704
rect 0 306008 800 306128
rect 356778 303560 357578 303680
rect 0 298120 800 298240
rect 356778 295536 357578 295656
rect 0 290232 800 290352
rect 356778 287512 357578 287632
rect 0 282344 800 282464
rect 356778 279488 357578 279608
rect 0 274456 800 274576
rect 356778 271464 357578 271584
rect 0 266568 800 266688
rect 356778 263440 357578 263560
rect 0 258680 800 258800
rect 356778 255416 357578 255536
rect 0 250792 800 250912
rect 356778 247392 357578 247512
rect 0 242904 800 243024
rect 356778 239368 357578 239488
rect 0 235016 800 235136
rect 356778 231344 357578 231464
rect 0 227128 800 227248
rect 356778 223320 357578 223440
rect 0 219240 800 219360
rect 356778 215296 357578 215416
rect 0 211352 800 211472
rect 356778 207272 357578 207392
rect 0 203464 800 203584
rect 356778 199248 357578 199368
rect 0 195576 800 195696
rect 356778 191224 357578 191344
rect 0 187688 800 187808
rect 356778 183200 357578 183320
rect 0 179800 800 179920
rect 356778 175176 357578 175296
rect 0 171912 800 172032
rect 356778 167152 357578 167272
rect 0 164024 800 164144
rect 356778 159128 357578 159248
rect 0 156136 800 156256
rect 356778 151104 357578 151224
rect 0 148248 800 148368
rect 356778 143080 357578 143200
rect 0 140360 800 140480
rect 356778 135056 357578 135176
rect 0 132472 800 132592
rect 356778 127032 357578 127152
rect 0 124584 800 124704
rect 356778 119008 357578 119128
rect 0 116696 800 116816
rect 356778 110984 357578 111104
rect 0 108808 800 108928
rect 356778 102960 357578 103080
rect 0 100920 800 101040
rect 356778 94936 357578 95056
rect 0 93032 800 93152
rect 356778 86912 357578 87032
rect 0 85144 800 85264
rect 356778 78888 357578 79008
rect 0 77256 800 77376
rect 356778 70864 357578 70984
rect 0 69368 800 69488
rect 356778 62840 357578 62960
rect 0 61480 800 61600
rect 356778 54816 357578 54936
rect 0 53592 800 53712
rect 356778 46792 357578 46912
rect 0 45704 800 45824
rect 356778 38768 357578 38888
rect 0 37816 800 37936
rect 356778 30744 357578 30864
rect 0 29928 800 30048
rect 356778 22720 357578 22840
rect 0 22040 800 22160
rect 356778 14696 357578 14816
rect 0 14152 800 14272
rect 356778 6672 357578 6792
rect 0 6264 800 6384
<< obsm3 >>
rect 800 424528 357090 428501
rect 880 424248 357090 424528
rect 800 424120 357090 424248
rect 800 423840 356698 424120
rect 800 416640 357090 423840
rect 880 416360 357090 416640
rect 800 416096 357090 416360
rect 800 415816 356698 416096
rect 800 408752 357090 415816
rect 880 408472 357090 408752
rect 800 408072 357090 408472
rect 800 407792 356698 408072
rect 800 400864 357090 407792
rect 880 400584 357090 400864
rect 800 400048 357090 400584
rect 800 399768 356698 400048
rect 800 392976 357090 399768
rect 880 392696 357090 392976
rect 800 392024 357090 392696
rect 800 391744 356698 392024
rect 800 385088 357090 391744
rect 880 384808 357090 385088
rect 800 384000 357090 384808
rect 800 383720 356698 384000
rect 800 377200 357090 383720
rect 880 376920 357090 377200
rect 800 375976 357090 376920
rect 800 375696 356698 375976
rect 800 369312 357090 375696
rect 880 369032 357090 369312
rect 800 367952 357090 369032
rect 800 367672 356698 367952
rect 800 361424 357090 367672
rect 880 361144 357090 361424
rect 800 359928 357090 361144
rect 800 359648 356698 359928
rect 800 353536 357090 359648
rect 880 353256 357090 353536
rect 800 351904 357090 353256
rect 800 351624 356698 351904
rect 800 345648 357090 351624
rect 880 345368 357090 345648
rect 800 343880 357090 345368
rect 800 343600 356698 343880
rect 800 337760 357090 343600
rect 880 337480 357090 337760
rect 800 335856 357090 337480
rect 800 335576 356698 335856
rect 800 329872 357090 335576
rect 880 329592 357090 329872
rect 800 327832 357090 329592
rect 800 327552 356698 327832
rect 800 321984 357090 327552
rect 880 321704 357090 321984
rect 800 319808 357090 321704
rect 800 319528 356698 319808
rect 800 314096 357090 319528
rect 880 313816 357090 314096
rect 800 311784 357090 313816
rect 800 311504 356698 311784
rect 800 306208 357090 311504
rect 880 305928 357090 306208
rect 800 303760 357090 305928
rect 800 303480 356698 303760
rect 800 298320 357090 303480
rect 880 298040 357090 298320
rect 800 295736 357090 298040
rect 800 295456 356698 295736
rect 800 290432 357090 295456
rect 880 290152 357090 290432
rect 800 287712 357090 290152
rect 800 287432 356698 287712
rect 800 282544 357090 287432
rect 880 282264 357090 282544
rect 800 279688 357090 282264
rect 800 279408 356698 279688
rect 800 274656 357090 279408
rect 880 274376 357090 274656
rect 800 271664 357090 274376
rect 800 271384 356698 271664
rect 800 266768 357090 271384
rect 880 266488 357090 266768
rect 800 263640 357090 266488
rect 800 263360 356698 263640
rect 800 258880 357090 263360
rect 880 258600 357090 258880
rect 800 255616 357090 258600
rect 800 255336 356698 255616
rect 800 250992 357090 255336
rect 880 250712 357090 250992
rect 800 247592 357090 250712
rect 800 247312 356698 247592
rect 800 243104 357090 247312
rect 880 242824 357090 243104
rect 800 239568 357090 242824
rect 800 239288 356698 239568
rect 800 235216 357090 239288
rect 880 234936 357090 235216
rect 800 231544 357090 234936
rect 800 231264 356698 231544
rect 800 227328 357090 231264
rect 880 227048 357090 227328
rect 800 223520 357090 227048
rect 800 223240 356698 223520
rect 800 219440 357090 223240
rect 880 219160 357090 219440
rect 800 215496 357090 219160
rect 800 215216 356698 215496
rect 800 211552 357090 215216
rect 880 211272 357090 211552
rect 800 207472 357090 211272
rect 800 207192 356698 207472
rect 800 203664 357090 207192
rect 880 203384 357090 203664
rect 800 199448 357090 203384
rect 800 199168 356698 199448
rect 800 195776 357090 199168
rect 880 195496 357090 195776
rect 800 191424 357090 195496
rect 800 191144 356698 191424
rect 800 187888 357090 191144
rect 880 187608 357090 187888
rect 800 183400 357090 187608
rect 800 183120 356698 183400
rect 800 180000 357090 183120
rect 880 179720 357090 180000
rect 800 175376 357090 179720
rect 800 175096 356698 175376
rect 800 172112 357090 175096
rect 880 171832 357090 172112
rect 800 167352 357090 171832
rect 800 167072 356698 167352
rect 800 164224 357090 167072
rect 880 163944 357090 164224
rect 800 159328 357090 163944
rect 800 159048 356698 159328
rect 800 156336 357090 159048
rect 880 156056 357090 156336
rect 800 151304 357090 156056
rect 800 151024 356698 151304
rect 800 148448 357090 151024
rect 880 148168 357090 148448
rect 800 143280 357090 148168
rect 800 143000 356698 143280
rect 800 140560 357090 143000
rect 880 140280 357090 140560
rect 800 135256 357090 140280
rect 800 134976 356698 135256
rect 800 132672 357090 134976
rect 880 132392 357090 132672
rect 800 127232 357090 132392
rect 800 126952 356698 127232
rect 800 124784 357090 126952
rect 880 124504 357090 124784
rect 800 119208 357090 124504
rect 800 118928 356698 119208
rect 800 116896 357090 118928
rect 880 116616 357090 116896
rect 800 111184 357090 116616
rect 800 110904 356698 111184
rect 800 109008 357090 110904
rect 880 108728 357090 109008
rect 800 103160 357090 108728
rect 800 102880 356698 103160
rect 800 101120 357090 102880
rect 880 100840 357090 101120
rect 800 95136 357090 100840
rect 800 94856 356698 95136
rect 800 93232 357090 94856
rect 880 92952 357090 93232
rect 800 87112 357090 92952
rect 800 86832 356698 87112
rect 800 85344 357090 86832
rect 880 85064 357090 85344
rect 800 79088 357090 85064
rect 800 78808 356698 79088
rect 800 77456 357090 78808
rect 880 77176 357090 77456
rect 800 71064 357090 77176
rect 800 70784 356698 71064
rect 800 69568 357090 70784
rect 880 69288 357090 69568
rect 800 63040 357090 69288
rect 800 62760 356698 63040
rect 800 61680 357090 62760
rect 880 61400 357090 61680
rect 800 55016 357090 61400
rect 800 54736 356698 55016
rect 800 53792 357090 54736
rect 880 53512 357090 53792
rect 800 46992 357090 53512
rect 800 46712 356698 46992
rect 800 45904 357090 46712
rect 880 45624 357090 45904
rect 800 38968 357090 45624
rect 800 38688 356698 38968
rect 800 38016 357090 38688
rect 880 37736 357090 38016
rect 800 30944 357090 37736
rect 800 30664 356698 30944
rect 800 30128 357090 30664
rect 880 29848 357090 30128
rect 800 22920 357090 29848
rect 800 22640 356698 22920
rect 800 22240 357090 22640
rect 880 21960 357090 22240
rect 800 14896 357090 21960
rect 800 14616 356698 14896
rect 800 14352 357090 14616
rect 880 14072 357090 14352
rect 800 6872 357090 14072
rect 800 6592 356698 6872
rect 800 6464 357090 6592
rect 880 6184 357090 6464
rect 800 2143 357090 6184
<< metal4 >>
rect 4208 2128 4528 428176
rect 19568 2128 19888 428176
rect 34928 2128 35248 428176
rect 50288 2128 50608 428176
rect 65648 2128 65968 428176
rect 81008 2128 81328 428176
rect 96368 2128 96688 428176
rect 111728 2128 112048 428176
rect 127088 2128 127408 428176
rect 142448 2128 142768 428176
rect 157808 2128 158128 428176
rect 173168 2128 173488 428176
rect 188528 2128 188848 428176
rect 203888 2128 204208 428176
rect 219248 2128 219568 428176
rect 234608 2128 234928 428176
rect 249968 2128 250288 428176
rect 265328 2128 265648 428176
rect 280688 2128 281008 428176
rect 296048 2128 296368 428176
rect 311408 2128 311728 428176
rect 326768 2128 327088 428176
rect 342128 2128 342448 428176
<< obsm4 >>
rect 1163 428256 357085 428501
rect 1163 3435 4128 428256
rect 4608 3435 19488 428256
rect 19968 3435 34848 428256
rect 35328 3435 50208 428256
rect 50688 3435 65568 428256
rect 66048 3435 80928 428256
rect 81408 3435 96288 428256
rect 96768 3435 111648 428256
rect 112128 3435 127008 428256
rect 127488 3435 142368 428256
rect 142848 3435 157728 428256
rect 158208 3435 173088 428256
rect 173568 3435 188448 428256
rect 188928 3435 203808 428256
rect 204288 3435 219168 428256
rect 219648 3435 234528 428256
rect 235008 3435 249888 428256
rect 250368 3435 265248 428256
rect 265728 3435 280608 428256
rect 281088 3435 295968 428256
rect 296448 3435 311328 428256
rect 311808 3435 326688 428256
rect 327168 3435 342048 428256
rect 342528 3435 357085 428256
<< labels >>
rlabel metal3 s 356778 175176 357578 175296 6 analog_io[0]
port 1 nsew signal bidirectional
rlabel metal2 s 272246 429996 272302 430796 6 analog_io[10]
port 2 nsew signal bidirectional
rlabel metal2 s 232870 429996 232926 430796 6 analog_io[11]
port 3 nsew signal bidirectional
rlabel metal2 s 193494 429996 193550 430796 6 analog_io[12]
port 4 nsew signal bidirectional
rlabel metal2 s 154118 429996 154174 430796 6 analog_io[13]
port 5 nsew signal bidirectional
rlabel metal2 s 114742 429996 114798 430796 6 analog_io[14]
port 6 nsew signal bidirectional
rlabel metal2 s 75366 429996 75422 430796 6 analog_io[15]
port 7 nsew signal bidirectional
rlabel metal2 s 35990 429996 36046 430796 6 analog_io[16]
port 8 nsew signal bidirectional
rlabel metal3 s 0 424328 800 424448 6 analog_io[17]
port 9 nsew signal bidirectional
rlabel metal3 s 0 392776 800 392896 6 analog_io[18]
port 10 nsew signal bidirectional
rlabel metal3 s 0 361224 800 361344 6 analog_io[19]
port 11 nsew signal bidirectional
rlabel metal3 s 356778 207272 357578 207392 6 analog_io[1]
port 12 nsew signal bidirectional
rlabel metal3 s 0 329672 800 329792 6 analog_io[20]
port 13 nsew signal bidirectional
rlabel metal3 s 0 298120 800 298240 6 analog_io[21]
port 14 nsew signal bidirectional
rlabel metal3 s 0 266568 800 266688 6 analog_io[22]
port 15 nsew signal bidirectional
rlabel metal3 s 0 235016 800 235136 6 analog_io[23]
port 16 nsew signal bidirectional
rlabel metal3 s 0 203464 800 203584 6 analog_io[24]
port 17 nsew signal bidirectional
rlabel metal3 s 0 171912 800 172032 6 analog_io[25]
port 18 nsew signal bidirectional
rlabel metal3 s 0 140360 800 140480 6 analog_io[26]
port 19 nsew signal bidirectional
rlabel metal3 s 0 108808 800 108928 6 analog_io[27]
port 20 nsew signal bidirectional
rlabel metal3 s 0 77256 800 77376 6 analog_io[28]
port 21 nsew signal bidirectional
rlabel metal3 s 356778 239368 357578 239488 6 analog_io[2]
port 22 nsew signal bidirectional
rlabel metal3 s 356778 271464 357578 271584 6 analog_io[3]
port 23 nsew signal bidirectional
rlabel metal3 s 356778 303560 357578 303680 6 analog_io[4]
port 24 nsew signal bidirectional
rlabel metal3 s 356778 335656 357578 335776 6 analog_io[5]
port 25 nsew signal bidirectional
rlabel metal3 s 356778 367752 357578 367872 6 analog_io[6]
port 26 nsew signal bidirectional
rlabel metal3 s 356778 399848 357578 399968 6 analog_io[7]
port 27 nsew signal bidirectional
rlabel metal2 s 350998 429996 351054 430796 6 analog_io[8]
port 28 nsew signal bidirectional
rlabel metal2 s 311622 429996 311678 430796 6 analog_io[9]
port 29 nsew signal bidirectional
rlabel metal3 s 356778 6672 357578 6792 6 io_in[0]
port 30 nsew signal input
rlabel metal3 s 356778 279488 357578 279608 6 io_in[10]
port 31 nsew signal input
rlabel metal3 s 356778 311584 357578 311704 6 io_in[11]
port 32 nsew signal input
rlabel metal3 s 356778 343680 357578 343800 6 io_in[12]
port 33 nsew signal input
rlabel metal3 s 356778 375776 357578 375896 6 io_in[13]
port 34 nsew signal input
rlabel metal3 s 356778 407872 357578 407992 6 io_in[14]
port 35 nsew signal input
rlabel metal2 s 341154 429996 341210 430796 6 io_in[15]
port 36 nsew signal input
rlabel metal2 s 301778 429996 301834 430796 6 io_in[16]
port 37 nsew signal input
rlabel metal2 s 262402 429996 262458 430796 6 io_in[17]
port 38 nsew signal input
rlabel metal2 s 223026 429996 223082 430796 6 io_in[18]
port 39 nsew signal input
rlabel metal2 s 183650 429996 183706 430796 6 io_in[19]
port 40 nsew signal input
rlabel metal3 s 356778 30744 357578 30864 6 io_in[1]
port 41 nsew signal input
rlabel metal2 s 144274 429996 144330 430796 6 io_in[20]
port 42 nsew signal input
rlabel metal2 s 104898 429996 104954 430796 6 io_in[21]
port 43 nsew signal input
rlabel metal2 s 65522 429996 65578 430796 6 io_in[22]
port 44 nsew signal input
rlabel metal2 s 26146 429996 26202 430796 6 io_in[23]
port 45 nsew signal input
rlabel metal3 s 0 416440 800 416560 6 io_in[24]
port 46 nsew signal input
rlabel metal3 s 0 384888 800 385008 6 io_in[25]
port 47 nsew signal input
rlabel metal3 s 0 353336 800 353456 6 io_in[26]
port 48 nsew signal input
rlabel metal3 s 0 321784 800 321904 6 io_in[27]
port 49 nsew signal input
rlabel metal3 s 0 290232 800 290352 6 io_in[28]
port 50 nsew signal input
rlabel metal3 s 0 258680 800 258800 6 io_in[29]
port 51 nsew signal input
rlabel metal3 s 356778 54816 357578 54936 6 io_in[2]
port 52 nsew signal input
rlabel metal3 s 0 227128 800 227248 6 io_in[30]
port 53 nsew signal input
rlabel metal3 s 0 195576 800 195696 6 io_in[31]
port 54 nsew signal input
rlabel metal3 s 0 164024 800 164144 6 io_in[32]
port 55 nsew signal input
rlabel metal3 s 0 132472 800 132592 6 io_in[33]
port 56 nsew signal input
rlabel metal3 s 0 100920 800 101040 6 io_in[34]
port 57 nsew signal input
rlabel metal3 s 0 69368 800 69488 6 io_in[35]
port 58 nsew signal input
rlabel metal3 s 0 45704 800 45824 6 io_in[36]
port 59 nsew signal input
rlabel metal3 s 0 22040 800 22160 6 io_in[37]
port 60 nsew signal input
rlabel metal3 s 356778 78888 357578 79008 6 io_in[3]
port 61 nsew signal input
rlabel metal3 s 356778 102960 357578 103080 6 io_in[4]
port 62 nsew signal input
rlabel metal3 s 356778 127032 357578 127152 6 io_in[5]
port 63 nsew signal input
rlabel metal3 s 356778 151104 357578 151224 6 io_in[6]
port 64 nsew signal input
rlabel metal3 s 356778 183200 357578 183320 6 io_in[7]
port 65 nsew signal input
rlabel metal3 s 356778 215296 357578 215416 6 io_in[8]
port 66 nsew signal input
rlabel metal3 s 356778 247392 357578 247512 6 io_in[9]
port 67 nsew signal input
rlabel metal3 s 356778 22720 357578 22840 6 io_oeb[0]
port 68 nsew signal output
rlabel metal3 s 356778 295536 357578 295656 6 io_oeb[10]
port 69 nsew signal output
rlabel metal3 s 356778 327632 357578 327752 6 io_oeb[11]
port 70 nsew signal output
rlabel metal3 s 356778 359728 357578 359848 6 io_oeb[12]
port 71 nsew signal output
rlabel metal3 s 356778 391824 357578 391944 6 io_oeb[13]
port 72 nsew signal output
rlabel metal3 s 356778 423920 357578 424040 6 io_oeb[14]
port 73 nsew signal output
rlabel metal2 s 321466 429996 321522 430796 6 io_oeb[15]
port 74 nsew signal output
rlabel metal2 s 282090 429996 282146 430796 6 io_oeb[16]
port 75 nsew signal output
rlabel metal2 s 242714 429996 242770 430796 6 io_oeb[17]
port 76 nsew signal output
rlabel metal2 s 203338 429996 203394 430796 6 io_oeb[18]
port 77 nsew signal output
rlabel metal2 s 163962 429996 164018 430796 6 io_oeb[19]
port 78 nsew signal output
rlabel metal3 s 356778 46792 357578 46912 6 io_oeb[1]
port 79 nsew signal output
rlabel metal2 s 124586 429996 124642 430796 6 io_oeb[20]
port 80 nsew signal output
rlabel metal2 s 85210 429996 85266 430796 6 io_oeb[21]
port 81 nsew signal output
rlabel metal2 s 45834 429996 45890 430796 6 io_oeb[22]
port 82 nsew signal output
rlabel metal2 s 6458 429996 6514 430796 6 io_oeb[23]
port 83 nsew signal output
rlabel metal3 s 0 400664 800 400784 6 io_oeb[24]
port 84 nsew signal output
rlabel metal3 s 0 369112 800 369232 6 io_oeb[25]
port 85 nsew signal output
rlabel metal3 s 0 337560 800 337680 6 io_oeb[26]
port 86 nsew signal output
rlabel metal3 s 0 306008 800 306128 6 io_oeb[27]
port 87 nsew signal output
rlabel metal3 s 0 274456 800 274576 6 io_oeb[28]
port 88 nsew signal output
rlabel metal3 s 0 242904 800 243024 6 io_oeb[29]
port 89 nsew signal output
rlabel metal3 s 356778 70864 357578 70984 6 io_oeb[2]
port 90 nsew signal output
rlabel metal3 s 0 211352 800 211472 6 io_oeb[30]
port 91 nsew signal output
rlabel metal3 s 0 179800 800 179920 6 io_oeb[31]
port 92 nsew signal output
rlabel metal3 s 0 148248 800 148368 6 io_oeb[32]
port 93 nsew signal output
rlabel metal3 s 0 116696 800 116816 6 io_oeb[33]
port 94 nsew signal output
rlabel metal3 s 0 85144 800 85264 6 io_oeb[34]
port 95 nsew signal output
rlabel metal3 s 0 53592 800 53712 6 io_oeb[35]
port 96 nsew signal output
rlabel metal3 s 0 29928 800 30048 6 io_oeb[36]
port 97 nsew signal output
rlabel metal3 s 0 6264 800 6384 6 io_oeb[37]
port 98 nsew signal output
rlabel metal3 s 356778 94936 357578 95056 6 io_oeb[3]
port 99 nsew signal output
rlabel metal3 s 356778 119008 357578 119128 6 io_oeb[4]
port 100 nsew signal output
rlabel metal3 s 356778 143080 357578 143200 6 io_oeb[5]
port 101 nsew signal output
rlabel metal3 s 356778 167152 357578 167272 6 io_oeb[6]
port 102 nsew signal output
rlabel metal3 s 356778 199248 357578 199368 6 io_oeb[7]
port 103 nsew signal output
rlabel metal3 s 356778 231344 357578 231464 6 io_oeb[8]
port 104 nsew signal output
rlabel metal3 s 356778 263440 357578 263560 6 io_oeb[9]
port 105 nsew signal output
rlabel metal3 s 356778 14696 357578 14816 6 io_out[0]
port 106 nsew signal output
rlabel metal3 s 356778 287512 357578 287632 6 io_out[10]
port 107 nsew signal output
rlabel metal3 s 356778 319608 357578 319728 6 io_out[11]
port 108 nsew signal output
rlabel metal3 s 356778 351704 357578 351824 6 io_out[12]
port 109 nsew signal output
rlabel metal3 s 356778 383800 357578 383920 6 io_out[13]
port 110 nsew signal output
rlabel metal3 s 356778 415896 357578 416016 6 io_out[14]
port 111 nsew signal output
rlabel metal2 s 331310 429996 331366 430796 6 io_out[15]
port 112 nsew signal output
rlabel metal2 s 291934 429996 291990 430796 6 io_out[16]
port 113 nsew signal output
rlabel metal2 s 252558 429996 252614 430796 6 io_out[17]
port 114 nsew signal output
rlabel metal2 s 213182 429996 213238 430796 6 io_out[18]
port 115 nsew signal output
rlabel metal2 s 173806 429996 173862 430796 6 io_out[19]
port 116 nsew signal output
rlabel metal3 s 356778 38768 357578 38888 6 io_out[1]
port 117 nsew signal output
rlabel metal2 s 134430 429996 134486 430796 6 io_out[20]
port 118 nsew signal output
rlabel metal2 s 95054 429996 95110 430796 6 io_out[21]
port 119 nsew signal output
rlabel metal2 s 55678 429996 55734 430796 6 io_out[22]
port 120 nsew signal output
rlabel metal2 s 16302 429996 16358 430796 6 io_out[23]
port 121 nsew signal output
rlabel metal3 s 0 408552 800 408672 6 io_out[24]
port 122 nsew signal output
rlabel metal3 s 0 377000 800 377120 6 io_out[25]
port 123 nsew signal output
rlabel metal3 s 0 345448 800 345568 6 io_out[26]
port 124 nsew signal output
rlabel metal3 s 0 313896 800 314016 6 io_out[27]
port 125 nsew signal output
rlabel metal3 s 0 282344 800 282464 6 io_out[28]
port 126 nsew signal output
rlabel metal3 s 0 250792 800 250912 6 io_out[29]
port 127 nsew signal output
rlabel metal3 s 356778 62840 357578 62960 6 io_out[2]
port 128 nsew signal output
rlabel metal3 s 0 219240 800 219360 6 io_out[30]
port 129 nsew signal output
rlabel metal3 s 0 187688 800 187808 6 io_out[31]
port 130 nsew signal output
rlabel metal3 s 0 156136 800 156256 6 io_out[32]
port 131 nsew signal output
rlabel metal3 s 0 124584 800 124704 6 io_out[33]
port 132 nsew signal output
rlabel metal3 s 0 93032 800 93152 6 io_out[34]
port 133 nsew signal output
rlabel metal3 s 0 61480 800 61600 6 io_out[35]
port 134 nsew signal output
rlabel metal3 s 0 37816 800 37936 6 io_out[36]
port 135 nsew signal output
rlabel metal3 s 0 14152 800 14272 6 io_out[37]
port 136 nsew signal output
rlabel metal3 s 356778 86912 357578 87032 6 io_out[3]
port 137 nsew signal output
rlabel metal3 s 356778 110984 357578 111104 6 io_out[4]
port 138 nsew signal output
rlabel metal3 s 356778 135056 357578 135176 6 io_out[5]
port 139 nsew signal output
rlabel metal3 s 356778 159128 357578 159248 6 io_out[6]
port 140 nsew signal output
rlabel metal3 s 356778 191224 357578 191344 6 io_out[7]
port 141 nsew signal output
rlabel metal3 s 356778 223320 357578 223440 6 io_out[8]
port 142 nsew signal output
rlabel metal3 s 356778 255416 357578 255536 6 io_out[9]
port 143 nsew signal output
rlabel metal2 s 88246 0 88302 800 6 la_data_in[0]
port 144 nsew signal input
rlabel metal2 s 281446 0 281502 800 6 la_data_in[100]
port 145 nsew signal input
rlabel metal2 s 283378 0 283434 800 6 la_data_in[101]
port 146 nsew signal input
rlabel metal2 s 285310 0 285366 800 6 la_data_in[102]
port 147 nsew signal input
rlabel metal2 s 287242 0 287298 800 6 la_data_in[103]
port 148 nsew signal input
rlabel metal2 s 289174 0 289230 800 6 la_data_in[104]
port 149 nsew signal input
rlabel metal2 s 291106 0 291162 800 6 la_data_in[105]
port 150 nsew signal input
rlabel metal2 s 293038 0 293094 800 6 la_data_in[106]
port 151 nsew signal input
rlabel metal2 s 294970 0 295026 800 6 la_data_in[107]
port 152 nsew signal input
rlabel metal2 s 296902 0 296958 800 6 la_data_in[108]
port 153 nsew signal input
rlabel metal2 s 298834 0 298890 800 6 la_data_in[109]
port 154 nsew signal input
rlabel metal2 s 107566 0 107622 800 6 la_data_in[10]
port 155 nsew signal input
rlabel metal2 s 300766 0 300822 800 6 la_data_in[110]
port 156 nsew signal input
rlabel metal2 s 302698 0 302754 800 6 la_data_in[111]
port 157 nsew signal input
rlabel metal2 s 304630 0 304686 800 6 la_data_in[112]
port 158 nsew signal input
rlabel metal2 s 306562 0 306618 800 6 la_data_in[113]
port 159 nsew signal input
rlabel metal2 s 308494 0 308550 800 6 la_data_in[114]
port 160 nsew signal input
rlabel metal2 s 310426 0 310482 800 6 la_data_in[115]
port 161 nsew signal input
rlabel metal2 s 312358 0 312414 800 6 la_data_in[116]
port 162 nsew signal input
rlabel metal2 s 314290 0 314346 800 6 la_data_in[117]
port 163 nsew signal input
rlabel metal2 s 316222 0 316278 800 6 la_data_in[118]
port 164 nsew signal input
rlabel metal2 s 318154 0 318210 800 6 la_data_in[119]
port 165 nsew signal input
rlabel metal2 s 109498 0 109554 800 6 la_data_in[11]
port 166 nsew signal input
rlabel metal2 s 320086 0 320142 800 6 la_data_in[120]
port 167 nsew signal input
rlabel metal2 s 322018 0 322074 800 6 la_data_in[121]
port 168 nsew signal input
rlabel metal2 s 323950 0 324006 800 6 la_data_in[122]
port 169 nsew signal input
rlabel metal2 s 325882 0 325938 800 6 la_data_in[123]
port 170 nsew signal input
rlabel metal2 s 327814 0 327870 800 6 la_data_in[124]
port 171 nsew signal input
rlabel metal2 s 329746 0 329802 800 6 la_data_in[125]
port 172 nsew signal input
rlabel metal2 s 331678 0 331734 800 6 la_data_in[126]
port 173 nsew signal input
rlabel metal2 s 333610 0 333666 800 6 la_data_in[127]
port 174 nsew signal input
rlabel metal2 s 111430 0 111486 800 6 la_data_in[12]
port 175 nsew signal input
rlabel metal2 s 113362 0 113418 800 6 la_data_in[13]
port 176 nsew signal input
rlabel metal2 s 115294 0 115350 800 6 la_data_in[14]
port 177 nsew signal input
rlabel metal2 s 117226 0 117282 800 6 la_data_in[15]
port 178 nsew signal input
rlabel metal2 s 119158 0 119214 800 6 la_data_in[16]
port 179 nsew signal input
rlabel metal2 s 121090 0 121146 800 6 la_data_in[17]
port 180 nsew signal input
rlabel metal2 s 123022 0 123078 800 6 la_data_in[18]
port 181 nsew signal input
rlabel metal2 s 124954 0 125010 800 6 la_data_in[19]
port 182 nsew signal input
rlabel metal2 s 90178 0 90234 800 6 la_data_in[1]
port 183 nsew signal input
rlabel metal2 s 126886 0 126942 800 6 la_data_in[20]
port 184 nsew signal input
rlabel metal2 s 128818 0 128874 800 6 la_data_in[21]
port 185 nsew signal input
rlabel metal2 s 130750 0 130806 800 6 la_data_in[22]
port 186 nsew signal input
rlabel metal2 s 132682 0 132738 800 6 la_data_in[23]
port 187 nsew signal input
rlabel metal2 s 134614 0 134670 800 6 la_data_in[24]
port 188 nsew signal input
rlabel metal2 s 136546 0 136602 800 6 la_data_in[25]
port 189 nsew signal input
rlabel metal2 s 138478 0 138534 800 6 la_data_in[26]
port 190 nsew signal input
rlabel metal2 s 140410 0 140466 800 6 la_data_in[27]
port 191 nsew signal input
rlabel metal2 s 142342 0 142398 800 6 la_data_in[28]
port 192 nsew signal input
rlabel metal2 s 144274 0 144330 800 6 la_data_in[29]
port 193 nsew signal input
rlabel metal2 s 92110 0 92166 800 6 la_data_in[2]
port 194 nsew signal input
rlabel metal2 s 146206 0 146262 800 6 la_data_in[30]
port 195 nsew signal input
rlabel metal2 s 148138 0 148194 800 6 la_data_in[31]
port 196 nsew signal input
rlabel metal2 s 150070 0 150126 800 6 la_data_in[32]
port 197 nsew signal input
rlabel metal2 s 152002 0 152058 800 6 la_data_in[33]
port 198 nsew signal input
rlabel metal2 s 153934 0 153990 800 6 la_data_in[34]
port 199 nsew signal input
rlabel metal2 s 155866 0 155922 800 6 la_data_in[35]
port 200 nsew signal input
rlabel metal2 s 157798 0 157854 800 6 la_data_in[36]
port 201 nsew signal input
rlabel metal2 s 159730 0 159786 800 6 la_data_in[37]
port 202 nsew signal input
rlabel metal2 s 161662 0 161718 800 6 la_data_in[38]
port 203 nsew signal input
rlabel metal2 s 163594 0 163650 800 6 la_data_in[39]
port 204 nsew signal input
rlabel metal2 s 94042 0 94098 800 6 la_data_in[3]
port 205 nsew signal input
rlabel metal2 s 165526 0 165582 800 6 la_data_in[40]
port 206 nsew signal input
rlabel metal2 s 167458 0 167514 800 6 la_data_in[41]
port 207 nsew signal input
rlabel metal2 s 169390 0 169446 800 6 la_data_in[42]
port 208 nsew signal input
rlabel metal2 s 171322 0 171378 800 6 la_data_in[43]
port 209 nsew signal input
rlabel metal2 s 173254 0 173310 800 6 la_data_in[44]
port 210 nsew signal input
rlabel metal2 s 175186 0 175242 800 6 la_data_in[45]
port 211 nsew signal input
rlabel metal2 s 177118 0 177174 800 6 la_data_in[46]
port 212 nsew signal input
rlabel metal2 s 179050 0 179106 800 6 la_data_in[47]
port 213 nsew signal input
rlabel metal2 s 180982 0 181038 800 6 la_data_in[48]
port 214 nsew signal input
rlabel metal2 s 182914 0 182970 800 6 la_data_in[49]
port 215 nsew signal input
rlabel metal2 s 95974 0 96030 800 6 la_data_in[4]
port 216 nsew signal input
rlabel metal2 s 184846 0 184902 800 6 la_data_in[50]
port 217 nsew signal input
rlabel metal2 s 186778 0 186834 800 6 la_data_in[51]
port 218 nsew signal input
rlabel metal2 s 188710 0 188766 800 6 la_data_in[52]
port 219 nsew signal input
rlabel metal2 s 190642 0 190698 800 6 la_data_in[53]
port 220 nsew signal input
rlabel metal2 s 192574 0 192630 800 6 la_data_in[54]
port 221 nsew signal input
rlabel metal2 s 194506 0 194562 800 6 la_data_in[55]
port 222 nsew signal input
rlabel metal2 s 196438 0 196494 800 6 la_data_in[56]
port 223 nsew signal input
rlabel metal2 s 198370 0 198426 800 6 la_data_in[57]
port 224 nsew signal input
rlabel metal2 s 200302 0 200358 800 6 la_data_in[58]
port 225 nsew signal input
rlabel metal2 s 202234 0 202290 800 6 la_data_in[59]
port 226 nsew signal input
rlabel metal2 s 97906 0 97962 800 6 la_data_in[5]
port 227 nsew signal input
rlabel metal2 s 204166 0 204222 800 6 la_data_in[60]
port 228 nsew signal input
rlabel metal2 s 206098 0 206154 800 6 la_data_in[61]
port 229 nsew signal input
rlabel metal2 s 208030 0 208086 800 6 la_data_in[62]
port 230 nsew signal input
rlabel metal2 s 209962 0 210018 800 6 la_data_in[63]
port 231 nsew signal input
rlabel metal2 s 211894 0 211950 800 6 la_data_in[64]
port 232 nsew signal input
rlabel metal2 s 213826 0 213882 800 6 la_data_in[65]
port 233 nsew signal input
rlabel metal2 s 215758 0 215814 800 6 la_data_in[66]
port 234 nsew signal input
rlabel metal2 s 217690 0 217746 800 6 la_data_in[67]
port 235 nsew signal input
rlabel metal2 s 219622 0 219678 800 6 la_data_in[68]
port 236 nsew signal input
rlabel metal2 s 221554 0 221610 800 6 la_data_in[69]
port 237 nsew signal input
rlabel metal2 s 99838 0 99894 800 6 la_data_in[6]
port 238 nsew signal input
rlabel metal2 s 223486 0 223542 800 6 la_data_in[70]
port 239 nsew signal input
rlabel metal2 s 225418 0 225474 800 6 la_data_in[71]
port 240 nsew signal input
rlabel metal2 s 227350 0 227406 800 6 la_data_in[72]
port 241 nsew signal input
rlabel metal2 s 229282 0 229338 800 6 la_data_in[73]
port 242 nsew signal input
rlabel metal2 s 231214 0 231270 800 6 la_data_in[74]
port 243 nsew signal input
rlabel metal2 s 233146 0 233202 800 6 la_data_in[75]
port 244 nsew signal input
rlabel metal2 s 235078 0 235134 800 6 la_data_in[76]
port 245 nsew signal input
rlabel metal2 s 237010 0 237066 800 6 la_data_in[77]
port 246 nsew signal input
rlabel metal2 s 238942 0 238998 800 6 la_data_in[78]
port 247 nsew signal input
rlabel metal2 s 240874 0 240930 800 6 la_data_in[79]
port 248 nsew signal input
rlabel metal2 s 101770 0 101826 800 6 la_data_in[7]
port 249 nsew signal input
rlabel metal2 s 242806 0 242862 800 6 la_data_in[80]
port 250 nsew signal input
rlabel metal2 s 244738 0 244794 800 6 la_data_in[81]
port 251 nsew signal input
rlabel metal2 s 246670 0 246726 800 6 la_data_in[82]
port 252 nsew signal input
rlabel metal2 s 248602 0 248658 800 6 la_data_in[83]
port 253 nsew signal input
rlabel metal2 s 250534 0 250590 800 6 la_data_in[84]
port 254 nsew signal input
rlabel metal2 s 252466 0 252522 800 6 la_data_in[85]
port 255 nsew signal input
rlabel metal2 s 254398 0 254454 800 6 la_data_in[86]
port 256 nsew signal input
rlabel metal2 s 256330 0 256386 800 6 la_data_in[87]
port 257 nsew signal input
rlabel metal2 s 258262 0 258318 800 6 la_data_in[88]
port 258 nsew signal input
rlabel metal2 s 260194 0 260250 800 6 la_data_in[89]
port 259 nsew signal input
rlabel metal2 s 103702 0 103758 800 6 la_data_in[8]
port 260 nsew signal input
rlabel metal2 s 262126 0 262182 800 6 la_data_in[90]
port 261 nsew signal input
rlabel metal2 s 264058 0 264114 800 6 la_data_in[91]
port 262 nsew signal input
rlabel metal2 s 265990 0 266046 800 6 la_data_in[92]
port 263 nsew signal input
rlabel metal2 s 267922 0 267978 800 6 la_data_in[93]
port 264 nsew signal input
rlabel metal2 s 269854 0 269910 800 6 la_data_in[94]
port 265 nsew signal input
rlabel metal2 s 271786 0 271842 800 6 la_data_in[95]
port 266 nsew signal input
rlabel metal2 s 273718 0 273774 800 6 la_data_in[96]
port 267 nsew signal input
rlabel metal2 s 275650 0 275706 800 6 la_data_in[97]
port 268 nsew signal input
rlabel metal2 s 277582 0 277638 800 6 la_data_in[98]
port 269 nsew signal input
rlabel metal2 s 279514 0 279570 800 6 la_data_in[99]
port 270 nsew signal input
rlabel metal2 s 105634 0 105690 800 6 la_data_in[9]
port 271 nsew signal input
rlabel metal2 s 88890 0 88946 800 6 la_data_out[0]
port 272 nsew signal output
rlabel metal2 s 282090 0 282146 800 6 la_data_out[100]
port 273 nsew signal output
rlabel metal2 s 284022 0 284078 800 6 la_data_out[101]
port 274 nsew signal output
rlabel metal2 s 285954 0 286010 800 6 la_data_out[102]
port 275 nsew signal output
rlabel metal2 s 287886 0 287942 800 6 la_data_out[103]
port 276 nsew signal output
rlabel metal2 s 289818 0 289874 800 6 la_data_out[104]
port 277 nsew signal output
rlabel metal2 s 291750 0 291806 800 6 la_data_out[105]
port 278 nsew signal output
rlabel metal2 s 293682 0 293738 800 6 la_data_out[106]
port 279 nsew signal output
rlabel metal2 s 295614 0 295670 800 6 la_data_out[107]
port 280 nsew signal output
rlabel metal2 s 297546 0 297602 800 6 la_data_out[108]
port 281 nsew signal output
rlabel metal2 s 299478 0 299534 800 6 la_data_out[109]
port 282 nsew signal output
rlabel metal2 s 108210 0 108266 800 6 la_data_out[10]
port 283 nsew signal output
rlabel metal2 s 301410 0 301466 800 6 la_data_out[110]
port 284 nsew signal output
rlabel metal2 s 303342 0 303398 800 6 la_data_out[111]
port 285 nsew signal output
rlabel metal2 s 305274 0 305330 800 6 la_data_out[112]
port 286 nsew signal output
rlabel metal2 s 307206 0 307262 800 6 la_data_out[113]
port 287 nsew signal output
rlabel metal2 s 309138 0 309194 800 6 la_data_out[114]
port 288 nsew signal output
rlabel metal2 s 311070 0 311126 800 6 la_data_out[115]
port 289 nsew signal output
rlabel metal2 s 313002 0 313058 800 6 la_data_out[116]
port 290 nsew signal output
rlabel metal2 s 314934 0 314990 800 6 la_data_out[117]
port 291 nsew signal output
rlabel metal2 s 316866 0 316922 800 6 la_data_out[118]
port 292 nsew signal output
rlabel metal2 s 318798 0 318854 800 6 la_data_out[119]
port 293 nsew signal output
rlabel metal2 s 110142 0 110198 800 6 la_data_out[11]
port 294 nsew signal output
rlabel metal2 s 320730 0 320786 800 6 la_data_out[120]
port 295 nsew signal output
rlabel metal2 s 322662 0 322718 800 6 la_data_out[121]
port 296 nsew signal output
rlabel metal2 s 324594 0 324650 800 6 la_data_out[122]
port 297 nsew signal output
rlabel metal2 s 326526 0 326582 800 6 la_data_out[123]
port 298 nsew signal output
rlabel metal2 s 328458 0 328514 800 6 la_data_out[124]
port 299 nsew signal output
rlabel metal2 s 330390 0 330446 800 6 la_data_out[125]
port 300 nsew signal output
rlabel metal2 s 332322 0 332378 800 6 la_data_out[126]
port 301 nsew signal output
rlabel metal2 s 334254 0 334310 800 6 la_data_out[127]
port 302 nsew signal output
rlabel metal2 s 112074 0 112130 800 6 la_data_out[12]
port 303 nsew signal output
rlabel metal2 s 114006 0 114062 800 6 la_data_out[13]
port 304 nsew signal output
rlabel metal2 s 115938 0 115994 800 6 la_data_out[14]
port 305 nsew signal output
rlabel metal2 s 117870 0 117926 800 6 la_data_out[15]
port 306 nsew signal output
rlabel metal2 s 119802 0 119858 800 6 la_data_out[16]
port 307 nsew signal output
rlabel metal2 s 121734 0 121790 800 6 la_data_out[17]
port 308 nsew signal output
rlabel metal2 s 123666 0 123722 800 6 la_data_out[18]
port 309 nsew signal output
rlabel metal2 s 125598 0 125654 800 6 la_data_out[19]
port 310 nsew signal output
rlabel metal2 s 90822 0 90878 800 6 la_data_out[1]
port 311 nsew signal output
rlabel metal2 s 127530 0 127586 800 6 la_data_out[20]
port 312 nsew signal output
rlabel metal2 s 129462 0 129518 800 6 la_data_out[21]
port 313 nsew signal output
rlabel metal2 s 131394 0 131450 800 6 la_data_out[22]
port 314 nsew signal output
rlabel metal2 s 133326 0 133382 800 6 la_data_out[23]
port 315 nsew signal output
rlabel metal2 s 135258 0 135314 800 6 la_data_out[24]
port 316 nsew signal output
rlabel metal2 s 137190 0 137246 800 6 la_data_out[25]
port 317 nsew signal output
rlabel metal2 s 139122 0 139178 800 6 la_data_out[26]
port 318 nsew signal output
rlabel metal2 s 141054 0 141110 800 6 la_data_out[27]
port 319 nsew signal output
rlabel metal2 s 142986 0 143042 800 6 la_data_out[28]
port 320 nsew signal output
rlabel metal2 s 144918 0 144974 800 6 la_data_out[29]
port 321 nsew signal output
rlabel metal2 s 92754 0 92810 800 6 la_data_out[2]
port 322 nsew signal output
rlabel metal2 s 146850 0 146906 800 6 la_data_out[30]
port 323 nsew signal output
rlabel metal2 s 148782 0 148838 800 6 la_data_out[31]
port 324 nsew signal output
rlabel metal2 s 150714 0 150770 800 6 la_data_out[32]
port 325 nsew signal output
rlabel metal2 s 152646 0 152702 800 6 la_data_out[33]
port 326 nsew signal output
rlabel metal2 s 154578 0 154634 800 6 la_data_out[34]
port 327 nsew signal output
rlabel metal2 s 156510 0 156566 800 6 la_data_out[35]
port 328 nsew signal output
rlabel metal2 s 158442 0 158498 800 6 la_data_out[36]
port 329 nsew signal output
rlabel metal2 s 160374 0 160430 800 6 la_data_out[37]
port 330 nsew signal output
rlabel metal2 s 162306 0 162362 800 6 la_data_out[38]
port 331 nsew signal output
rlabel metal2 s 164238 0 164294 800 6 la_data_out[39]
port 332 nsew signal output
rlabel metal2 s 94686 0 94742 800 6 la_data_out[3]
port 333 nsew signal output
rlabel metal2 s 166170 0 166226 800 6 la_data_out[40]
port 334 nsew signal output
rlabel metal2 s 168102 0 168158 800 6 la_data_out[41]
port 335 nsew signal output
rlabel metal2 s 170034 0 170090 800 6 la_data_out[42]
port 336 nsew signal output
rlabel metal2 s 171966 0 172022 800 6 la_data_out[43]
port 337 nsew signal output
rlabel metal2 s 173898 0 173954 800 6 la_data_out[44]
port 338 nsew signal output
rlabel metal2 s 175830 0 175886 800 6 la_data_out[45]
port 339 nsew signal output
rlabel metal2 s 177762 0 177818 800 6 la_data_out[46]
port 340 nsew signal output
rlabel metal2 s 179694 0 179750 800 6 la_data_out[47]
port 341 nsew signal output
rlabel metal2 s 181626 0 181682 800 6 la_data_out[48]
port 342 nsew signal output
rlabel metal2 s 183558 0 183614 800 6 la_data_out[49]
port 343 nsew signal output
rlabel metal2 s 96618 0 96674 800 6 la_data_out[4]
port 344 nsew signal output
rlabel metal2 s 185490 0 185546 800 6 la_data_out[50]
port 345 nsew signal output
rlabel metal2 s 187422 0 187478 800 6 la_data_out[51]
port 346 nsew signal output
rlabel metal2 s 189354 0 189410 800 6 la_data_out[52]
port 347 nsew signal output
rlabel metal2 s 191286 0 191342 800 6 la_data_out[53]
port 348 nsew signal output
rlabel metal2 s 193218 0 193274 800 6 la_data_out[54]
port 349 nsew signal output
rlabel metal2 s 195150 0 195206 800 6 la_data_out[55]
port 350 nsew signal output
rlabel metal2 s 197082 0 197138 800 6 la_data_out[56]
port 351 nsew signal output
rlabel metal2 s 199014 0 199070 800 6 la_data_out[57]
port 352 nsew signal output
rlabel metal2 s 200946 0 201002 800 6 la_data_out[58]
port 353 nsew signal output
rlabel metal2 s 202878 0 202934 800 6 la_data_out[59]
port 354 nsew signal output
rlabel metal2 s 98550 0 98606 800 6 la_data_out[5]
port 355 nsew signal output
rlabel metal2 s 204810 0 204866 800 6 la_data_out[60]
port 356 nsew signal output
rlabel metal2 s 206742 0 206798 800 6 la_data_out[61]
port 357 nsew signal output
rlabel metal2 s 208674 0 208730 800 6 la_data_out[62]
port 358 nsew signal output
rlabel metal2 s 210606 0 210662 800 6 la_data_out[63]
port 359 nsew signal output
rlabel metal2 s 212538 0 212594 800 6 la_data_out[64]
port 360 nsew signal output
rlabel metal2 s 214470 0 214526 800 6 la_data_out[65]
port 361 nsew signal output
rlabel metal2 s 216402 0 216458 800 6 la_data_out[66]
port 362 nsew signal output
rlabel metal2 s 218334 0 218390 800 6 la_data_out[67]
port 363 nsew signal output
rlabel metal2 s 220266 0 220322 800 6 la_data_out[68]
port 364 nsew signal output
rlabel metal2 s 222198 0 222254 800 6 la_data_out[69]
port 365 nsew signal output
rlabel metal2 s 100482 0 100538 800 6 la_data_out[6]
port 366 nsew signal output
rlabel metal2 s 224130 0 224186 800 6 la_data_out[70]
port 367 nsew signal output
rlabel metal2 s 226062 0 226118 800 6 la_data_out[71]
port 368 nsew signal output
rlabel metal2 s 227994 0 228050 800 6 la_data_out[72]
port 369 nsew signal output
rlabel metal2 s 229926 0 229982 800 6 la_data_out[73]
port 370 nsew signal output
rlabel metal2 s 231858 0 231914 800 6 la_data_out[74]
port 371 nsew signal output
rlabel metal2 s 233790 0 233846 800 6 la_data_out[75]
port 372 nsew signal output
rlabel metal2 s 235722 0 235778 800 6 la_data_out[76]
port 373 nsew signal output
rlabel metal2 s 237654 0 237710 800 6 la_data_out[77]
port 374 nsew signal output
rlabel metal2 s 239586 0 239642 800 6 la_data_out[78]
port 375 nsew signal output
rlabel metal2 s 241518 0 241574 800 6 la_data_out[79]
port 376 nsew signal output
rlabel metal2 s 102414 0 102470 800 6 la_data_out[7]
port 377 nsew signal output
rlabel metal2 s 243450 0 243506 800 6 la_data_out[80]
port 378 nsew signal output
rlabel metal2 s 245382 0 245438 800 6 la_data_out[81]
port 379 nsew signal output
rlabel metal2 s 247314 0 247370 800 6 la_data_out[82]
port 380 nsew signal output
rlabel metal2 s 249246 0 249302 800 6 la_data_out[83]
port 381 nsew signal output
rlabel metal2 s 251178 0 251234 800 6 la_data_out[84]
port 382 nsew signal output
rlabel metal2 s 253110 0 253166 800 6 la_data_out[85]
port 383 nsew signal output
rlabel metal2 s 255042 0 255098 800 6 la_data_out[86]
port 384 nsew signal output
rlabel metal2 s 256974 0 257030 800 6 la_data_out[87]
port 385 nsew signal output
rlabel metal2 s 258906 0 258962 800 6 la_data_out[88]
port 386 nsew signal output
rlabel metal2 s 260838 0 260894 800 6 la_data_out[89]
port 387 nsew signal output
rlabel metal2 s 104346 0 104402 800 6 la_data_out[8]
port 388 nsew signal output
rlabel metal2 s 262770 0 262826 800 6 la_data_out[90]
port 389 nsew signal output
rlabel metal2 s 264702 0 264758 800 6 la_data_out[91]
port 390 nsew signal output
rlabel metal2 s 266634 0 266690 800 6 la_data_out[92]
port 391 nsew signal output
rlabel metal2 s 268566 0 268622 800 6 la_data_out[93]
port 392 nsew signal output
rlabel metal2 s 270498 0 270554 800 6 la_data_out[94]
port 393 nsew signal output
rlabel metal2 s 272430 0 272486 800 6 la_data_out[95]
port 394 nsew signal output
rlabel metal2 s 274362 0 274418 800 6 la_data_out[96]
port 395 nsew signal output
rlabel metal2 s 276294 0 276350 800 6 la_data_out[97]
port 396 nsew signal output
rlabel metal2 s 278226 0 278282 800 6 la_data_out[98]
port 397 nsew signal output
rlabel metal2 s 280158 0 280214 800 6 la_data_out[99]
port 398 nsew signal output
rlabel metal2 s 106278 0 106334 800 6 la_data_out[9]
port 399 nsew signal output
rlabel metal2 s 89534 0 89590 800 6 la_oenb[0]
port 400 nsew signal input
rlabel metal2 s 282734 0 282790 800 6 la_oenb[100]
port 401 nsew signal input
rlabel metal2 s 284666 0 284722 800 6 la_oenb[101]
port 402 nsew signal input
rlabel metal2 s 286598 0 286654 800 6 la_oenb[102]
port 403 nsew signal input
rlabel metal2 s 288530 0 288586 800 6 la_oenb[103]
port 404 nsew signal input
rlabel metal2 s 290462 0 290518 800 6 la_oenb[104]
port 405 nsew signal input
rlabel metal2 s 292394 0 292450 800 6 la_oenb[105]
port 406 nsew signal input
rlabel metal2 s 294326 0 294382 800 6 la_oenb[106]
port 407 nsew signal input
rlabel metal2 s 296258 0 296314 800 6 la_oenb[107]
port 408 nsew signal input
rlabel metal2 s 298190 0 298246 800 6 la_oenb[108]
port 409 nsew signal input
rlabel metal2 s 300122 0 300178 800 6 la_oenb[109]
port 410 nsew signal input
rlabel metal2 s 108854 0 108910 800 6 la_oenb[10]
port 411 nsew signal input
rlabel metal2 s 302054 0 302110 800 6 la_oenb[110]
port 412 nsew signal input
rlabel metal2 s 303986 0 304042 800 6 la_oenb[111]
port 413 nsew signal input
rlabel metal2 s 305918 0 305974 800 6 la_oenb[112]
port 414 nsew signal input
rlabel metal2 s 307850 0 307906 800 6 la_oenb[113]
port 415 nsew signal input
rlabel metal2 s 309782 0 309838 800 6 la_oenb[114]
port 416 nsew signal input
rlabel metal2 s 311714 0 311770 800 6 la_oenb[115]
port 417 nsew signal input
rlabel metal2 s 313646 0 313702 800 6 la_oenb[116]
port 418 nsew signal input
rlabel metal2 s 315578 0 315634 800 6 la_oenb[117]
port 419 nsew signal input
rlabel metal2 s 317510 0 317566 800 6 la_oenb[118]
port 420 nsew signal input
rlabel metal2 s 319442 0 319498 800 6 la_oenb[119]
port 421 nsew signal input
rlabel metal2 s 110786 0 110842 800 6 la_oenb[11]
port 422 nsew signal input
rlabel metal2 s 321374 0 321430 800 6 la_oenb[120]
port 423 nsew signal input
rlabel metal2 s 323306 0 323362 800 6 la_oenb[121]
port 424 nsew signal input
rlabel metal2 s 325238 0 325294 800 6 la_oenb[122]
port 425 nsew signal input
rlabel metal2 s 327170 0 327226 800 6 la_oenb[123]
port 426 nsew signal input
rlabel metal2 s 329102 0 329158 800 6 la_oenb[124]
port 427 nsew signal input
rlabel metal2 s 331034 0 331090 800 6 la_oenb[125]
port 428 nsew signal input
rlabel metal2 s 332966 0 333022 800 6 la_oenb[126]
port 429 nsew signal input
rlabel metal2 s 334898 0 334954 800 6 la_oenb[127]
port 430 nsew signal input
rlabel metal2 s 112718 0 112774 800 6 la_oenb[12]
port 431 nsew signal input
rlabel metal2 s 114650 0 114706 800 6 la_oenb[13]
port 432 nsew signal input
rlabel metal2 s 116582 0 116638 800 6 la_oenb[14]
port 433 nsew signal input
rlabel metal2 s 118514 0 118570 800 6 la_oenb[15]
port 434 nsew signal input
rlabel metal2 s 120446 0 120502 800 6 la_oenb[16]
port 435 nsew signal input
rlabel metal2 s 122378 0 122434 800 6 la_oenb[17]
port 436 nsew signal input
rlabel metal2 s 124310 0 124366 800 6 la_oenb[18]
port 437 nsew signal input
rlabel metal2 s 126242 0 126298 800 6 la_oenb[19]
port 438 nsew signal input
rlabel metal2 s 91466 0 91522 800 6 la_oenb[1]
port 439 nsew signal input
rlabel metal2 s 128174 0 128230 800 6 la_oenb[20]
port 440 nsew signal input
rlabel metal2 s 130106 0 130162 800 6 la_oenb[21]
port 441 nsew signal input
rlabel metal2 s 132038 0 132094 800 6 la_oenb[22]
port 442 nsew signal input
rlabel metal2 s 133970 0 134026 800 6 la_oenb[23]
port 443 nsew signal input
rlabel metal2 s 135902 0 135958 800 6 la_oenb[24]
port 444 nsew signal input
rlabel metal2 s 137834 0 137890 800 6 la_oenb[25]
port 445 nsew signal input
rlabel metal2 s 139766 0 139822 800 6 la_oenb[26]
port 446 nsew signal input
rlabel metal2 s 141698 0 141754 800 6 la_oenb[27]
port 447 nsew signal input
rlabel metal2 s 143630 0 143686 800 6 la_oenb[28]
port 448 nsew signal input
rlabel metal2 s 145562 0 145618 800 6 la_oenb[29]
port 449 nsew signal input
rlabel metal2 s 93398 0 93454 800 6 la_oenb[2]
port 450 nsew signal input
rlabel metal2 s 147494 0 147550 800 6 la_oenb[30]
port 451 nsew signal input
rlabel metal2 s 149426 0 149482 800 6 la_oenb[31]
port 452 nsew signal input
rlabel metal2 s 151358 0 151414 800 6 la_oenb[32]
port 453 nsew signal input
rlabel metal2 s 153290 0 153346 800 6 la_oenb[33]
port 454 nsew signal input
rlabel metal2 s 155222 0 155278 800 6 la_oenb[34]
port 455 nsew signal input
rlabel metal2 s 157154 0 157210 800 6 la_oenb[35]
port 456 nsew signal input
rlabel metal2 s 159086 0 159142 800 6 la_oenb[36]
port 457 nsew signal input
rlabel metal2 s 161018 0 161074 800 6 la_oenb[37]
port 458 nsew signal input
rlabel metal2 s 162950 0 163006 800 6 la_oenb[38]
port 459 nsew signal input
rlabel metal2 s 164882 0 164938 800 6 la_oenb[39]
port 460 nsew signal input
rlabel metal2 s 95330 0 95386 800 6 la_oenb[3]
port 461 nsew signal input
rlabel metal2 s 166814 0 166870 800 6 la_oenb[40]
port 462 nsew signal input
rlabel metal2 s 168746 0 168802 800 6 la_oenb[41]
port 463 nsew signal input
rlabel metal2 s 170678 0 170734 800 6 la_oenb[42]
port 464 nsew signal input
rlabel metal2 s 172610 0 172666 800 6 la_oenb[43]
port 465 nsew signal input
rlabel metal2 s 174542 0 174598 800 6 la_oenb[44]
port 466 nsew signal input
rlabel metal2 s 176474 0 176530 800 6 la_oenb[45]
port 467 nsew signal input
rlabel metal2 s 178406 0 178462 800 6 la_oenb[46]
port 468 nsew signal input
rlabel metal2 s 180338 0 180394 800 6 la_oenb[47]
port 469 nsew signal input
rlabel metal2 s 182270 0 182326 800 6 la_oenb[48]
port 470 nsew signal input
rlabel metal2 s 184202 0 184258 800 6 la_oenb[49]
port 471 nsew signal input
rlabel metal2 s 97262 0 97318 800 6 la_oenb[4]
port 472 nsew signal input
rlabel metal2 s 186134 0 186190 800 6 la_oenb[50]
port 473 nsew signal input
rlabel metal2 s 188066 0 188122 800 6 la_oenb[51]
port 474 nsew signal input
rlabel metal2 s 189998 0 190054 800 6 la_oenb[52]
port 475 nsew signal input
rlabel metal2 s 191930 0 191986 800 6 la_oenb[53]
port 476 nsew signal input
rlabel metal2 s 193862 0 193918 800 6 la_oenb[54]
port 477 nsew signal input
rlabel metal2 s 195794 0 195850 800 6 la_oenb[55]
port 478 nsew signal input
rlabel metal2 s 197726 0 197782 800 6 la_oenb[56]
port 479 nsew signal input
rlabel metal2 s 199658 0 199714 800 6 la_oenb[57]
port 480 nsew signal input
rlabel metal2 s 201590 0 201646 800 6 la_oenb[58]
port 481 nsew signal input
rlabel metal2 s 203522 0 203578 800 6 la_oenb[59]
port 482 nsew signal input
rlabel metal2 s 99194 0 99250 800 6 la_oenb[5]
port 483 nsew signal input
rlabel metal2 s 205454 0 205510 800 6 la_oenb[60]
port 484 nsew signal input
rlabel metal2 s 207386 0 207442 800 6 la_oenb[61]
port 485 nsew signal input
rlabel metal2 s 209318 0 209374 800 6 la_oenb[62]
port 486 nsew signal input
rlabel metal2 s 211250 0 211306 800 6 la_oenb[63]
port 487 nsew signal input
rlabel metal2 s 213182 0 213238 800 6 la_oenb[64]
port 488 nsew signal input
rlabel metal2 s 215114 0 215170 800 6 la_oenb[65]
port 489 nsew signal input
rlabel metal2 s 217046 0 217102 800 6 la_oenb[66]
port 490 nsew signal input
rlabel metal2 s 218978 0 219034 800 6 la_oenb[67]
port 491 nsew signal input
rlabel metal2 s 220910 0 220966 800 6 la_oenb[68]
port 492 nsew signal input
rlabel metal2 s 222842 0 222898 800 6 la_oenb[69]
port 493 nsew signal input
rlabel metal2 s 101126 0 101182 800 6 la_oenb[6]
port 494 nsew signal input
rlabel metal2 s 224774 0 224830 800 6 la_oenb[70]
port 495 nsew signal input
rlabel metal2 s 226706 0 226762 800 6 la_oenb[71]
port 496 nsew signal input
rlabel metal2 s 228638 0 228694 800 6 la_oenb[72]
port 497 nsew signal input
rlabel metal2 s 230570 0 230626 800 6 la_oenb[73]
port 498 nsew signal input
rlabel metal2 s 232502 0 232558 800 6 la_oenb[74]
port 499 nsew signal input
rlabel metal2 s 234434 0 234490 800 6 la_oenb[75]
port 500 nsew signal input
rlabel metal2 s 236366 0 236422 800 6 la_oenb[76]
port 501 nsew signal input
rlabel metal2 s 238298 0 238354 800 6 la_oenb[77]
port 502 nsew signal input
rlabel metal2 s 240230 0 240286 800 6 la_oenb[78]
port 503 nsew signal input
rlabel metal2 s 242162 0 242218 800 6 la_oenb[79]
port 504 nsew signal input
rlabel metal2 s 103058 0 103114 800 6 la_oenb[7]
port 505 nsew signal input
rlabel metal2 s 244094 0 244150 800 6 la_oenb[80]
port 506 nsew signal input
rlabel metal2 s 246026 0 246082 800 6 la_oenb[81]
port 507 nsew signal input
rlabel metal2 s 247958 0 248014 800 6 la_oenb[82]
port 508 nsew signal input
rlabel metal2 s 249890 0 249946 800 6 la_oenb[83]
port 509 nsew signal input
rlabel metal2 s 251822 0 251878 800 6 la_oenb[84]
port 510 nsew signal input
rlabel metal2 s 253754 0 253810 800 6 la_oenb[85]
port 511 nsew signal input
rlabel metal2 s 255686 0 255742 800 6 la_oenb[86]
port 512 nsew signal input
rlabel metal2 s 257618 0 257674 800 6 la_oenb[87]
port 513 nsew signal input
rlabel metal2 s 259550 0 259606 800 6 la_oenb[88]
port 514 nsew signal input
rlabel metal2 s 261482 0 261538 800 6 la_oenb[89]
port 515 nsew signal input
rlabel metal2 s 104990 0 105046 800 6 la_oenb[8]
port 516 nsew signal input
rlabel metal2 s 263414 0 263470 800 6 la_oenb[90]
port 517 nsew signal input
rlabel metal2 s 265346 0 265402 800 6 la_oenb[91]
port 518 nsew signal input
rlabel metal2 s 267278 0 267334 800 6 la_oenb[92]
port 519 nsew signal input
rlabel metal2 s 269210 0 269266 800 6 la_oenb[93]
port 520 nsew signal input
rlabel metal2 s 271142 0 271198 800 6 la_oenb[94]
port 521 nsew signal input
rlabel metal2 s 273074 0 273130 800 6 la_oenb[95]
port 522 nsew signal input
rlabel metal2 s 275006 0 275062 800 6 la_oenb[96]
port 523 nsew signal input
rlabel metal2 s 276938 0 276994 800 6 la_oenb[97]
port 524 nsew signal input
rlabel metal2 s 278870 0 278926 800 6 la_oenb[98]
port 525 nsew signal input
rlabel metal2 s 280802 0 280858 800 6 la_oenb[99]
port 526 nsew signal input
rlabel metal2 s 106922 0 106978 800 6 la_oenb[9]
port 527 nsew signal input
rlabel metal2 s 335542 0 335598 800 6 user_clock2
port 528 nsew signal input
rlabel metal2 s 336186 0 336242 800 6 user_irq[0]
port 529 nsew signal output
rlabel metal2 s 336830 0 336886 800 6 user_irq[1]
port 530 nsew signal output
rlabel metal2 s 337474 0 337530 800 6 user_irq[2]
port 531 nsew signal output
rlabel metal4 s 4208 2128 4528 428176 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 428176 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 65648 2128 65968 428176 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 96368 2128 96688 428176 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 127088 2128 127408 428176 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 157808 2128 158128 428176 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 188528 2128 188848 428176 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 219248 2128 219568 428176 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 249968 2128 250288 428176 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 280688 2128 281008 428176 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 311408 2128 311728 428176 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 342128 2128 342448 428176 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 19568 2128 19888 428176 6 vssd1
port 533 nsew ground bidirectional
rlabel metal4 s 50288 2128 50608 428176 6 vssd1
port 533 nsew ground bidirectional
rlabel metal4 s 81008 2128 81328 428176 6 vssd1
port 533 nsew ground bidirectional
rlabel metal4 s 111728 2128 112048 428176 6 vssd1
port 533 nsew ground bidirectional
rlabel metal4 s 142448 2128 142768 428176 6 vssd1
port 533 nsew ground bidirectional
rlabel metal4 s 173168 2128 173488 428176 6 vssd1
port 533 nsew ground bidirectional
rlabel metal4 s 203888 2128 204208 428176 6 vssd1
port 533 nsew ground bidirectional
rlabel metal4 s 234608 2128 234928 428176 6 vssd1
port 533 nsew ground bidirectional
rlabel metal4 s 265328 2128 265648 428176 6 vssd1
port 533 nsew ground bidirectional
rlabel metal4 s 296048 2128 296368 428176 6 vssd1
port 533 nsew ground bidirectional
rlabel metal4 s 326768 2128 327088 428176 6 vssd1
port 533 nsew ground bidirectional
rlabel metal2 s 19982 0 20038 800 6 wb_clk_i
port 534 nsew signal input
rlabel metal2 s 20626 0 20682 800 6 wb_rst_i
port 535 nsew signal input
rlabel metal2 s 21270 0 21326 800 6 wbs_ack_o
port 536 nsew signal output
rlabel metal2 s 23846 0 23902 800 6 wbs_adr_i[0]
port 537 nsew signal input
rlabel metal2 s 45742 0 45798 800 6 wbs_adr_i[10]
port 538 nsew signal input
rlabel metal2 s 47674 0 47730 800 6 wbs_adr_i[11]
port 539 nsew signal input
rlabel metal2 s 49606 0 49662 800 6 wbs_adr_i[12]
port 540 nsew signal input
rlabel metal2 s 51538 0 51594 800 6 wbs_adr_i[13]
port 541 nsew signal input
rlabel metal2 s 53470 0 53526 800 6 wbs_adr_i[14]
port 542 nsew signal input
rlabel metal2 s 55402 0 55458 800 6 wbs_adr_i[15]
port 543 nsew signal input
rlabel metal2 s 57334 0 57390 800 6 wbs_adr_i[16]
port 544 nsew signal input
rlabel metal2 s 59266 0 59322 800 6 wbs_adr_i[17]
port 545 nsew signal input
rlabel metal2 s 61198 0 61254 800 6 wbs_adr_i[18]
port 546 nsew signal input
rlabel metal2 s 63130 0 63186 800 6 wbs_adr_i[19]
port 547 nsew signal input
rlabel metal2 s 26422 0 26478 800 6 wbs_adr_i[1]
port 548 nsew signal input
rlabel metal2 s 65062 0 65118 800 6 wbs_adr_i[20]
port 549 nsew signal input
rlabel metal2 s 66994 0 67050 800 6 wbs_adr_i[21]
port 550 nsew signal input
rlabel metal2 s 68926 0 68982 800 6 wbs_adr_i[22]
port 551 nsew signal input
rlabel metal2 s 70858 0 70914 800 6 wbs_adr_i[23]
port 552 nsew signal input
rlabel metal2 s 72790 0 72846 800 6 wbs_adr_i[24]
port 553 nsew signal input
rlabel metal2 s 74722 0 74778 800 6 wbs_adr_i[25]
port 554 nsew signal input
rlabel metal2 s 76654 0 76710 800 6 wbs_adr_i[26]
port 555 nsew signal input
rlabel metal2 s 78586 0 78642 800 6 wbs_adr_i[27]
port 556 nsew signal input
rlabel metal2 s 80518 0 80574 800 6 wbs_adr_i[28]
port 557 nsew signal input
rlabel metal2 s 82450 0 82506 800 6 wbs_adr_i[29]
port 558 nsew signal input
rlabel metal2 s 28998 0 29054 800 6 wbs_adr_i[2]
port 559 nsew signal input
rlabel metal2 s 84382 0 84438 800 6 wbs_adr_i[30]
port 560 nsew signal input
rlabel metal2 s 86314 0 86370 800 6 wbs_adr_i[31]
port 561 nsew signal input
rlabel metal2 s 31574 0 31630 800 6 wbs_adr_i[3]
port 562 nsew signal input
rlabel metal2 s 34150 0 34206 800 6 wbs_adr_i[4]
port 563 nsew signal input
rlabel metal2 s 36082 0 36138 800 6 wbs_adr_i[5]
port 564 nsew signal input
rlabel metal2 s 38014 0 38070 800 6 wbs_adr_i[6]
port 565 nsew signal input
rlabel metal2 s 39946 0 40002 800 6 wbs_adr_i[7]
port 566 nsew signal input
rlabel metal2 s 41878 0 41934 800 6 wbs_adr_i[8]
port 567 nsew signal input
rlabel metal2 s 43810 0 43866 800 6 wbs_adr_i[9]
port 568 nsew signal input
rlabel metal2 s 21914 0 21970 800 6 wbs_cyc_i
port 569 nsew signal input
rlabel metal2 s 24490 0 24546 800 6 wbs_dat_i[0]
port 570 nsew signal input
rlabel metal2 s 46386 0 46442 800 6 wbs_dat_i[10]
port 571 nsew signal input
rlabel metal2 s 48318 0 48374 800 6 wbs_dat_i[11]
port 572 nsew signal input
rlabel metal2 s 50250 0 50306 800 6 wbs_dat_i[12]
port 573 nsew signal input
rlabel metal2 s 52182 0 52238 800 6 wbs_dat_i[13]
port 574 nsew signal input
rlabel metal2 s 54114 0 54170 800 6 wbs_dat_i[14]
port 575 nsew signal input
rlabel metal2 s 56046 0 56102 800 6 wbs_dat_i[15]
port 576 nsew signal input
rlabel metal2 s 57978 0 58034 800 6 wbs_dat_i[16]
port 577 nsew signal input
rlabel metal2 s 59910 0 59966 800 6 wbs_dat_i[17]
port 578 nsew signal input
rlabel metal2 s 61842 0 61898 800 6 wbs_dat_i[18]
port 579 nsew signal input
rlabel metal2 s 63774 0 63830 800 6 wbs_dat_i[19]
port 580 nsew signal input
rlabel metal2 s 27066 0 27122 800 6 wbs_dat_i[1]
port 581 nsew signal input
rlabel metal2 s 65706 0 65762 800 6 wbs_dat_i[20]
port 582 nsew signal input
rlabel metal2 s 67638 0 67694 800 6 wbs_dat_i[21]
port 583 nsew signal input
rlabel metal2 s 69570 0 69626 800 6 wbs_dat_i[22]
port 584 nsew signal input
rlabel metal2 s 71502 0 71558 800 6 wbs_dat_i[23]
port 585 nsew signal input
rlabel metal2 s 73434 0 73490 800 6 wbs_dat_i[24]
port 586 nsew signal input
rlabel metal2 s 75366 0 75422 800 6 wbs_dat_i[25]
port 587 nsew signal input
rlabel metal2 s 77298 0 77354 800 6 wbs_dat_i[26]
port 588 nsew signal input
rlabel metal2 s 79230 0 79286 800 6 wbs_dat_i[27]
port 589 nsew signal input
rlabel metal2 s 81162 0 81218 800 6 wbs_dat_i[28]
port 590 nsew signal input
rlabel metal2 s 83094 0 83150 800 6 wbs_dat_i[29]
port 591 nsew signal input
rlabel metal2 s 29642 0 29698 800 6 wbs_dat_i[2]
port 592 nsew signal input
rlabel metal2 s 85026 0 85082 800 6 wbs_dat_i[30]
port 593 nsew signal input
rlabel metal2 s 86958 0 87014 800 6 wbs_dat_i[31]
port 594 nsew signal input
rlabel metal2 s 32218 0 32274 800 6 wbs_dat_i[3]
port 595 nsew signal input
rlabel metal2 s 34794 0 34850 800 6 wbs_dat_i[4]
port 596 nsew signal input
rlabel metal2 s 36726 0 36782 800 6 wbs_dat_i[5]
port 597 nsew signal input
rlabel metal2 s 38658 0 38714 800 6 wbs_dat_i[6]
port 598 nsew signal input
rlabel metal2 s 40590 0 40646 800 6 wbs_dat_i[7]
port 599 nsew signal input
rlabel metal2 s 42522 0 42578 800 6 wbs_dat_i[8]
port 600 nsew signal input
rlabel metal2 s 44454 0 44510 800 6 wbs_dat_i[9]
port 601 nsew signal input
rlabel metal2 s 25134 0 25190 800 6 wbs_dat_o[0]
port 602 nsew signal output
rlabel metal2 s 47030 0 47086 800 6 wbs_dat_o[10]
port 603 nsew signal output
rlabel metal2 s 48962 0 49018 800 6 wbs_dat_o[11]
port 604 nsew signal output
rlabel metal2 s 50894 0 50950 800 6 wbs_dat_o[12]
port 605 nsew signal output
rlabel metal2 s 52826 0 52882 800 6 wbs_dat_o[13]
port 606 nsew signal output
rlabel metal2 s 54758 0 54814 800 6 wbs_dat_o[14]
port 607 nsew signal output
rlabel metal2 s 56690 0 56746 800 6 wbs_dat_o[15]
port 608 nsew signal output
rlabel metal2 s 58622 0 58678 800 6 wbs_dat_o[16]
port 609 nsew signal output
rlabel metal2 s 60554 0 60610 800 6 wbs_dat_o[17]
port 610 nsew signal output
rlabel metal2 s 62486 0 62542 800 6 wbs_dat_o[18]
port 611 nsew signal output
rlabel metal2 s 64418 0 64474 800 6 wbs_dat_o[19]
port 612 nsew signal output
rlabel metal2 s 27710 0 27766 800 6 wbs_dat_o[1]
port 613 nsew signal output
rlabel metal2 s 66350 0 66406 800 6 wbs_dat_o[20]
port 614 nsew signal output
rlabel metal2 s 68282 0 68338 800 6 wbs_dat_o[21]
port 615 nsew signal output
rlabel metal2 s 70214 0 70270 800 6 wbs_dat_o[22]
port 616 nsew signal output
rlabel metal2 s 72146 0 72202 800 6 wbs_dat_o[23]
port 617 nsew signal output
rlabel metal2 s 74078 0 74134 800 6 wbs_dat_o[24]
port 618 nsew signal output
rlabel metal2 s 76010 0 76066 800 6 wbs_dat_o[25]
port 619 nsew signal output
rlabel metal2 s 77942 0 77998 800 6 wbs_dat_o[26]
port 620 nsew signal output
rlabel metal2 s 79874 0 79930 800 6 wbs_dat_o[27]
port 621 nsew signal output
rlabel metal2 s 81806 0 81862 800 6 wbs_dat_o[28]
port 622 nsew signal output
rlabel metal2 s 83738 0 83794 800 6 wbs_dat_o[29]
port 623 nsew signal output
rlabel metal2 s 30286 0 30342 800 6 wbs_dat_o[2]
port 624 nsew signal output
rlabel metal2 s 85670 0 85726 800 6 wbs_dat_o[30]
port 625 nsew signal output
rlabel metal2 s 87602 0 87658 800 6 wbs_dat_o[31]
port 626 nsew signal output
rlabel metal2 s 32862 0 32918 800 6 wbs_dat_o[3]
port 627 nsew signal output
rlabel metal2 s 35438 0 35494 800 6 wbs_dat_o[4]
port 628 nsew signal output
rlabel metal2 s 37370 0 37426 800 6 wbs_dat_o[5]
port 629 nsew signal output
rlabel metal2 s 39302 0 39358 800 6 wbs_dat_o[6]
port 630 nsew signal output
rlabel metal2 s 41234 0 41290 800 6 wbs_dat_o[7]
port 631 nsew signal output
rlabel metal2 s 43166 0 43222 800 6 wbs_dat_o[8]
port 632 nsew signal output
rlabel metal2 s 45098 0 45154 800 6 wbs_dat_o[9]
port 633 nsew signal output
rlabel metal2 s 25778 0 25834 800 6 wbs_sel_i[0]
port 634 nsew signal input
rlabel metal2 s 28354 0 28410 800 6 wbs_sel_i[1]
port 635 nsew signal input
rlabel metal2 s 30930 0 30986 800 6 wbs_sel_i[2]
port 636 nsew signal input
rlabel metal2 s 33506 0 33562 800 6 wbs_sel_i[3]
port 637 nsew signal input
rlabel metal2 s 22558 0 22614 800 6 wbs_stb_i
port 638 nsew signal input
rlabel metal2 s 23202 0 23258 800 6 wbs_we_i
port 639 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 357578 430796
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 346380922
string GDS_FILE /mnt/r/work/Rift2Go_2300_Sky130_MPW8/openlane/user_proj_example/runs/22_12_21_10_35/results/signoff/rift2Wrap.magic.gds
string GDS_START 1856444
<< end >>

